��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω������?9X�1�Z�U���T��ײ2��>���^k�/7�?1�(�c��ly[�$D֍C95^T��6\Xa��7��Į�N��=i�@x_\q[�@�0�I���j{�N<��;��� B]�pE���	x]̃Dj#^Da����M�[�.�sj��
�M��ļz����)�,�˛D��w���旴4�����:��@���b���$[G��m$�;�`��v��p�㈍x���t�켻�S���c,31�-elwB(�93;2���Zߧl4���0�?�1~�x�c�>j����d��S�W�>��Q�d����t�mR��:�����-��3���7�Jk�b#Ӡe��?�F��&��;�Éi���W:�*c��,v˶�9�ĒTC��0��`�R&.1� 0��]�������yW�u���;���A��j`��'�����`U+n%K)��k��Ǣ���N�y�Yc���;��sD���L�S5H�j.F�{��>�a��{��/Ƽ���\�4�s���rH
>TT	q��$�2�����b��ǾI}`�~�MUs �?oQ�%'�s����o���_�xm7��(С�"pX�����U�?��+�x�8�n����Oq:m�j�{_5Jwʛ���[E�8z���U ��?��k�Jd����r�>>7�*���/���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc������2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h~09h�i�Nq�{5��]�0�lK'���Xw����Q4?���ʢ\��|�����o�3ts�JFAa�ߖ�g��o�4��?����DNZ�j׫���?_W�\I��ఽ��`g�5��!08/?�s�m/C�N{a�9O!JoE'U�Y�y��
r�)�Y¹w����i��T!ix�AH�k[�^��_6�L�r��W�����%3?���kW���;��sD���L�S5H�j.F��%�	�r��L�Xڈ*-}|��ι%9��oGo�Z�J��ݪ�nX�#fZC��磋��w.V&��B֥�(����5���ռ�j��I���j{�܆L(,�Tf1}Kط��4q����S��Ǵ��BR�^Ƒ�ӥ�e%)>�Z��&��J�1�KB|1<\w¹��<d����n���u3v��U̢�Ab�%^T_.�z0"���	�9K��b?��]��E*�h3��{I�B�+�7m_T���Q��K���ma��y�~��ۢ>�xn^%��+0�l�R<�q��f�}���D)��!�`�(i3�o��C!T*Y�{'%s���'����F�r�f�t��6��	���`y������q��ww�=�J�5Y%T��BPS�)37J*uc�A�L'R�o�����5�%]���a(􆿳�ټ*w2�56�[b�0<��c��Et�Y�{'%s��.|Z���I7��-5��6��	���`y����ꢤ�Og�ś� ����]�!��	Ǹ�y85�����څ��;�¬pX��g��U-�eן�-�Q�Z�M��<��z��}�\w��0]�9+�����o��C!T*�q���U����?�N�By3��<Z鎬�����X���*_��(֥�S�)37J*u>����CΫa������<��z��}���w�V�"-4��h�]8+��T����oGo�Z�������--�p�,Xs1ܢzk˷NË�����8��z{��E�EYZ/�矘��-n��I�?g�f��Qө}�i���W:SJr���S =�M�ߚ�zy�g���+
���C�gAO��ً�}�Y�ןw�8���/����Z1`� k�|6�8>�
�����g�,P�n^P��:w�(�����@^7&ģM�)sWmyY��!둿8(?�3���Ib����rs�i�jf� l�Ǜ������CyW�f�tR�wX��}�
�?�k {P@2���4��)�ep�G;w�b!��u��5?�&P-�"z�a<�Y�{'%s���'����F�r�f�t��6��	���`y����@����gGT���/ ����C�#�,Z鎬�������(���P����ˮ��lC��U�T�\ ��i3�|)sՀ�T:���V���)(��8��d�٣��c�A�L'��!�a��5�%]���a(􆿳���2����.��DP֞ ?h�	9��v�n`5�fK��0z�cULjaGkƊ~F˯�+)�"j���b7���Øf�ƫ�G���N���T	6:��=����זρ5�D��
∺V��܅t�iZ]XF�������́&�Ө��{�V�f��[��iJ�~�Y���(���;����f!�`�(i3�i3<�f�D���X���`>����������o��)�ak�m6"�,�>E��ʆ�In��tT?�7G|`���N�v*$�!�`�(i3�i3<�f�D���X���`����"��5�w�yzw�����+"�,�>E��4];ˍH��!�,���;���2[����|��1�J�a3mPy�S�W�W`!�`�(i3x�]�V���t�����[F�a�+S:H��+܆"BT�(��c����L�{7�ܥ��2�`e7��9��×�>�濖��#�(y"BT�(��c����L�{���D	��U�l>o��|���bǬ�= �zbw��(2�����
�b��{�P}�=]A��O�T=�4e=��-Y�VN�=���Ζ�{QU2����0�5tU���+�J��U<o^.K�}/��<Ӭ�/�"�����_G��?u:�L��Y%T��BP��&��J�UG�s����s�٩���I���Т��^�\7�ܥ��2�`e7��9���I^Ɍ؝�hy�/B/���^!l���Z1����x�'aU<o^.K�}qW8+���?iRPs�&�Ө��{�}+�o�n��iJ�~�Y���(��U��?D��!�`�(i3"�,�>E��ʆ�In��tT?�7G|`~�Y���(�M����H}R!�`�(i3"�,�>E��ʆ�In��tT?�7G|`���N���96!�`�(i3"�,�>E��ʆ�In��t�_�R�Gl�����b���V�Lx{<qH�~�"�,�>E��4];ˍH��\B�����g�q~[{Q�|�\m��Z��N�l�B�r���E����F���8�TPm=_g}b��t�S:H��+܆��K����!�`�(i3зq8�Ј)w�<�_N�-Ł$��Ь>�#�_���}Dq�f��.��Ԕ�]��3a��!�`�(i3���D	��U�l>o��|���bǬ�=l�����2�����
����7
"�,�>E��4];ˍH����TI��Ԫ,щ�"�t� ��O���}���i!�`�(i3���+�J��U<o^.K�}�d	c�b��8���&�r��SQQv�x�����D ML:��Yg6���=�4e=��-"w߻Y��}Dq�f�(����O�^�|n�M�!�`�(i3���D	��U�l>o��|���JLm|��|#HK��@=���b�A������!�`�(i37�ܥ��2�`e7��9��×�>���`�)J*~���f�A�������E����F���8�TP��@E�`�8���&�'�al��pz!�
�W@!�`�(i3=]A��O�T=�4e=��-Y�VN�=���Ζ�{QU2���A������!�`�(i3x�]�V���t�����[F�a�+#�n�%�<�'`ٲ�,�Xʚ@hY%T��BP��&��J�UG�s����s�٩���I����:�Y���зq8�Ј)w�<�_NX�ʟ�3���M&������h�? "a��%}w�dN����+�J��U<o^.K�}qW8+����8���&����uSj��Q�s΁�a�n��=]A��O�T=�4e=��-��~��A��<�6�Q=	�H�Z����Q��nT��Q#>[��b�-W��^[�΍�>!�`�(i3!�`�(i3���+�J��U<o^.K�}5��s� �+U���z�W�F��X�C+�t̷@V�� �!�`�(i3!�`�(i3Y%T��BP��&��J����$�!h�SSB�����m�%��~?H�?���i�jw�jս�������8�TP��k��p�ݹ��}��Z&�lq6�.ʲPdLG���6!�`�(i3!�`�(i37�ܥ��2����*����i��>�`vx��c6�����b(!�`�(i3!�`�(i3"�,�>E��4];ˍH�v��K.Ū�X��oҍvx��c6������|)i��OP���!�`�(i3"�,�>E��4];ˍH�v��K.Ū�X��oҍ�`��rE����ij~�*k`Ë��!�`�(i3"�,�>E��ʆ�In��t�_�R�G��!=.�
kZ)� [��v���Q:�g�a2�-�!�`�(i3x�]�V��w�7qyX����1��H,\ͨ܉p������aUMf�n�Q]�����	!�`�(i37�ܥ��2��fƆ���?|5#�Gm�X:��+��N�C��(4];ˍH�T֟��B�:УWKŃ
.�Ūz�ȣ)[CȪ�U� ���_��z���u�;����2e�5�O֐V���o��k�I#�ā9���8����W�%kԒ�P�K�T�b��M��d��p∺V��܅\4L$ֵ�j�iy[���ҋX����Q��C� ��!�`�(i3!�`�(i3!�`�(i3k��j �%��:wJ~��b{'�t���s�����s|Nb��'1-��B�Noq�ށ �~K[���#<��z��}�z�-~BLI�!�`�(i3!�`�(i3!�`�(i3V����(��N!��qő��{����gFUӮY�E��vNd�)i���
�mN�By3��<Z鎬����a�gN�3c!�`�(i3!�`�(i3!�`�(i3�����U�#�ҒIs{��f��C�'��"�����q��l0q�\E��0j�iy[���ҋX������S8�=	���/lg������T�\ ���KD��}[e��0�U�S{����<�6�Q=$�D5�bY[XҹvXI)�vNd�)i+�0\�NN�By3��<Z鎬�������(���$�~����$^�V]��}1;Z�减l|�*"k���(ӈ��4��S;UA7��I+N����-���q\��Zt%��m&<g+b󆤐=��{l�f|��rs�i���YN�聟�lҟ�,0=]^	�&|#9���� л�.���N���>���n�J�LQ��w�6�5�p����}���S�)37J*uc�A�L'�t�O5u�l�+�	�g��U-�ee�@Rv����my$�N��;� ��b�� л�o���ߞ����>���n
�z��+?i`YS���*';���3�q���Um��#��*y��+�^@��#	Ͼ7�Z#^L�)�4)	���E7��I+��v��q��y�&؏R!׻�p���f
�@"��wҦ�kQW֑��bk<����-�˳k�L��<�6�Q=�w�3����f
�@"��g�����Mgs�4�����DW+'4"��.B�2g>~qA��@����M�P�;�ȓM�Me���섫�So#ȓM�Me��x�2�Hxl�� ޘ_�9��\�'�������>Q��?qr��Kl3��T�Ҹ�MS�B�|��T��tn�+�e��j�3����&Y��V�贅����OD��G͘B./�<ĩ�46�;:���t�b|bQ��� Ǐ˨�g���!G#�<��z��}�<ͧ�:|�"��ӌ�r,�ttT� O���hZ鎬����=���ޒC>ž_�F���^W��kD���4B'�e��n�FM��`��\n$̱~"��>d�c#�'����^W��k�������!�`�(i3!�`�(i3�Ѳ��aS�!-�+_����1�"`��Ę*��7��S��>z��OP�/#�x�+-�+q�!�`�(i3!�`�(i3i`YS�����9Z������?6z�9�ot8��$��.A��+��T��s�٩��um8:8���]�!��5��E0����|e"� 䉇o�M���!O@T'���Xw�����U�VA�ڦ�c4&bݷ�%O�e��n00�8��P6�Y��\���(����A-u��6�0;��ȓM�Me����ΜtȓM�Me��x�2�Hxl�� ޘ_�9��\�'�U�"�����<º#xH�i�é���Vs��nlH�I<�6�Q=�w�3����f
�@"��g�����R��H�O��	�d[��K�pHj�4�\��F���77AƐ^�87��I+�T���B�H��y�&؏R!׻�p���f
�@"tL�^VG����L1�%TԞ}�{J��n��&�P��k<kbm�ѕ����[�|�"u��ӳ��C1��g��U��q�o�u�/ZB�JU��\bE����Kl3��+�I,�S���R����)�&��_���c�.DٖM?�_�9���{l�f|��:2QYeƈ)P<�ܓ�Y竷b��"&�����'�Z鎬����Ĺ#{��ž_�Fȓ'�al��p�M>�I�dB��{l�f|��:2QYeƈ)P<�ܓ�YSƏw0���:ʽ�f0�J.�A�]�!���\B��Vƺ'���g�>k0�ޏ�OEǄ���]�!��	Ǹ�y85��q幊s�?����H�n�f���\�g��U-�ee�@Rv����my$�N��;� ��b�� л���eY�b6=,����hQ���}Q'݀�=��⹌y��o��C!T*Y�{'%sgeߪ�{$�~����$�⹌y�S�UE^����Cҷ��e�ˇ�h����2�[Q	��
�Q�}#�ҒIs{S�>��{A��"�����f��z�� л��Ujc(h�t�%ho����G���r(�:�f,��iQ��e�Z鎬�������(����} "m��^�V]��}Г����ѓ�1���`���A�O
i�c�r׶|�ل�\I��w��,c�A�L'�t�O#��XvU(�8���/�7��I+�:����fSM0.��4;�. ��F����U�e	�K~9M=�6��#eCL�x��m��58*������,��ٙ���O�Dw
�
�{��_r�e~5�O�%E#P�⒍~��$�x�Wt!�`�(i3!�`�(i3!�`�(i3J�a$�Y  �VBD�!��"��{�R�ܯ	�J3��Iћ<��!�`�(i3!�`�(i3!�`�(i3Ǒ�e}5��Ь��z�q�\E��0���/�!�`�(i3!�`�(i3!�`�(i3!�`�(i3v{��lw	~�'�eo�ANL�P����<����t�T�V�r��}�������y�:Fa�7����Q+��
ņANL��ʡ.>��5�5���/9�=eSe.��a��o���H�RtV�^�� ߌ��!�`�(i3!�`�(i3!�`�(i3!�`�(i3?��ِ���I��<��;b�-�2��;�P�t�5W?�;�끷�Q+��
ņANL�P����<��m)�X�\
<�7�C��!�`�(i3�U��)���yk;�C>��ӚH�RtV�^�璓�c�������t �[l;M?��y�!�`�(i3G��ô��b���0��!�`�(i3!�`�(i3!�`�(i3.�T�w��'�i�*ڶ�UKs,��(��{�Oh0����v�9���+��9,(W ���t�1tSjv�V�Ո����oz�N۞��n�!�`�(i3�uz�#-]ix��?�S��h0�����1�>`�nT���t!h�ݚ�Н����F��O��;b�-�2��;�P�t�5W?�;���z��O�&�Z�%�k�.�g3Z�j5�{�CL�x��m_�/��!N\PPE�H�b"�uQ��z/�B{�o
�s��$�Z;��|B[g�� ���S�@�
37�˱�5PM�^-q�x�l��1:�N�*�x��0�C�D^J����'�kf�<�IUR5�(<�%by&6����u*_g5��pC50
���=:�<��W{0`�ǣ©����8���w�������K�7����;�줦�ݚ�Н��zsO%!E���tR�/p.0��I�![�Do�9�ݚ�Н�d�hb{;!�`�(i3���u�UgF˯�+)��&�C�/:��+���y��̨X&|a�#�I7��-5��5Z��¥�����-��+�&-��A�sxW�O�,��L���D:����ЊQvN�G!�`�(i3B�O�%J(V�K=�u��!�`�(i3�.E�f\���dv��oTN֢&@��&�MQNv�2���w0��U젩`#�4>?� �1SƏw0��-��2Q��	3H����'���Xw�j�7��j�n�y�f�?ǉ�=J�a3mPy�x�6�
Xg�%Y��̗0z�cUL0:_\�c��,5�)�F�B�'��a�U�xn�Oq-����b=���hy��:�KZ����b=���hy�_�⥳�"_�X;p`�YmC,iguY��j3������i�b{����"�2��}��g��9|P�X;p`���C�,�4��؟O�,�Xʚ@h-��?�l�`��!�`�(i3�57�0q��&8�,��A��=5<�!�d�<�.�g3Z�j5�{���������Rr������ ���D�]Z�Vy}'��vr��-��2.[��9�GͿK�mJ�0�6�ETk/�0��nz�������b�G��S��e�Ul�;p�����4A���8�4%��0/3S��n��@IE�U����S8��y�)xʔ���V�� �\�HP@�a�;�k�fՂ��!O@T'���Xw%��[z����&4}��X�ҋX����7�8������q?����OEǄ���]�!��	Ǹ�y85��3}�@�7��?E/6Ұ��8_�|#9���jC�p���G�݈,��S�)37J*uc�A�L'����f�.`�G](p���*R�wX���d��<���])���/�Z鎬����a3sĹb��B���7{�ҋX������S8��y�)xʔ���V�� ���`y�����G���Ld�-P�Z:����"� X$L��~��0���u���xf36�x8@�*�p�q�BZS[]N���B
�����xf36�x8@�*�p�ɹ��I�N���B
�����xf36k""��{��P*N�2���2���n��y�5`P�~�v�r��Rϻt<� ).�x6��l���{Ф�E�+��c�4];ˍH���@E�`���f^��iT�v���5��L�����;�줦�ݚ�Н��|r��n����q��3[�W�W��<��W{0`�R����2�n���\��BO&j0��.@.?E��TZ����>�SS�]si�O�����rRV��F��s-"&`���*1�mJ�0�6��M��yr&VxI	��m+)q�����B�N��Q�>σwE����4���"5���q�؅��FJ��/��<Ӭ�d�6��*@j ���N�����yc�b1���4];ˍH�m=_g}b��7ݲ����F!�f�t�x��~:@@!~�X����Ѵ���(�V*�u���1��؅��FJ��u6Mn+J�h�����mf_N2�CD�� ]IzL͊�q��C(�W�Ηfl��緺4v�r��Rϻx�]�V��v��K.Ū(T����ɻt��o�5������b7�ܥ��2�/��:M/�ա�^�jjl��緺4c�b1���4];ˍH�m=_g}b��7ݲ������勤U�@k����c�Zw|�pMGD@�F��qX�ʟ�H�Ѱ,���e���}����� NM�P����؅��FJ��qW8+����PK�k�V�t(]�XS����ڸłv#���ޑ؅��FJ��qW8+����PK�k�V�t(]�XS����ڸ��P����؅��FJ��qW8+������f^�	�q{dNJR�)��<|��}R�ElGD@�F��qW��Ґ�Yj:{b6��P'�gY%w�!,q��%�
��4];ˍH�T֟��BXaFg�N��%`���g�E�so��!�`�(i3u7btc�(ӫ�)F�9!�`�(i3!�`�(i3=]A��O�T=�4e=��-)����%�KW℀4��>ll��4?��X9���		���@!�`�(i3!�`�(i3JHn��z��r9�3k��u��aV$n������x���!�`�(i3!�`�(i3�E����F�'n�^0om�i�K�~sȸ�"rR�ԌY&�xL��$J��!�`�(i3!�`�(i3 ���3�ҺIÙ=�H���mL�02Y��kک��d��G�P�x�!�`�(i3!�`�(i3���D	��U�l>o��|���JLm|��� �5�v�l[��:���}M,�d��ҥ3�k�`�H��A������V�Ϯ4];ˍH�'N2��D����&�Q�,;#L�ܽU���¥������c�4��s���rۺ�!�`�(i3!�`�(i3JHn��z���G7��k��u��:��+���f�.`�Gy��̨!�`�(i3�E����F�'n�^0o�C�~��j��mJ�0�6�p)�?�{�7