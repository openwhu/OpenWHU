module AD_Data
(
	CLK, RSTn, AD_DigData_In, AD_CSn, AD_Clk, AD_Address, Data_Out, CS_Valid_Sig
);

	 input CLK;
	 input RSTn;		//SW0
	 
	 input AD_DigData_In;	 
	 output AD_CSn;
	 output AD_Clk;
	 output AD_Address;
	
	 output [9:0]Data_Out;	
	 output reg CS_Valid_Sig;
	 
	 reg AD_CSn_r;
	 reg AD_Clk_r;
	 reg AD_Address_r;
	 reg [9:0]Data_Out_r;
	 		 
     wire [3:0]Addr = 4'b0101;	   	//AIN5   
	 /*wire [3:0]Addr = 4'b1101;			//Verf+   */
	 /*wire [3:0]Addr = 4'b1011;			//（Verf+ + Verf-）/2*/
	 
/****************************************/		 
	 reg [7:0]Cnt1;
	 reg Cnt1_en;
	 
	always @ ( posedge CLK or negedge RSTn )
		begin
			if( !RSTn )
				begin
					Cnt1 <= 8'd0;
				end
			else if( Cnt1 == 8'd12 )						// generate " I/O CLOCK ( AD_Clk ) " , period is 2*13*20ns = 520ns
				begin
					Cnt1 <= 8'b0;
				end
			else if( Cnt1_en )
				begin
					Cnt1 <= Cnt1 + 1'b1;
				end
			else 
				Cnt1 <= 8'b0;			
		end

/****************************************/		
	 reg [7:0]Cnt2;
	 reg Cnt2_en;
	 
	always @ ( posedge CLK or negedge RSTn )
		begin
			if( !RSTn )
				begin
					Cnt2 <= 8'd0;
				end
		 	else if( Cnt2 == 8'd71 )		// generate " tsu(cs) " , Delayed Time is 72*20ns = 1440ns > 1.425us
				begin
					Cnt2 <= 8'b0;
				end 
			else if( Cnt2_en )
				begin
					Cnt2 <= Cnt2 + 1'b1;
				end
			else 
				Cnt2 <= 8'b0;			
		end
	
/********************************************/	
	 reg [7:0]Cnt3;
	 reg Cnt3_en;

	always @ ( posedge CLK or negedge RSTn )
		begin
			if( !RSTn )
				begin
					Cnt3 <= 8'd0;
				end
		 	else if( Cnt3 == 8'd25 )		// generate a clock signal to control the data transmitted to "AD_Address", 													
				begin								//	period is 26*20ns = 520ns			
					Cnt3 <= 8'b0;
				end 
			else if( Cnt3_en )
				begin
					Cnt3 <= Cnt3 + 1'b1;
				end
			else 
				Cnt3 <= 8'b0;			
		end	
	
/*****************************************/	
	 reg [10:0]Cnt4;
	 reg Cnt4_en;

	always @ ( posedge CLK or negedge RSTn )
		begin
			if( !RSTn )
				begin
					Cnt4 <= 11'd0;
				end
		 	else if( Cnt4 == 11'd1050 )		// generate " Conversion time " , Delayed Time is 1050*20ns = 21us
				begin								 
					Cnt4 <= 11'b0;	
				end 
			else if( Cnt4_en )
				begin
					Cnt4 <= Cnt4 + 1'b1;
				end
			else 
				Cnt4 <= 11'b0;			
		end
		
/*******************************************/	
	 reg [4:0]i;
	 
	always @ ( posedge CLK or negedge RSTn )
		begin
			if( !RSTn )
				begin
					i <= 5'b1;
					Data_Out_r <= 10'b0;					
					Cnt1_en <= 1'b0;
					Cnt2_en <= 1'b0;
					Cnt3_en <= 1'b0;
					Cnt4_en <= 1'b0;
					CS_Valid_Sig <= 1'b1;
				end
			else  	
				case( i )
					'd1: begin							//initial state
							AD_CSn_r <= 1'b1;
							AD_Clk_r <= 1'b0;
							Cnt1_en <= 1'b0;
							Cnt2_en <= 1'b0;
							Cnt3_en <= 1'b0;
							Cnt4_en <= 1'b0;
							i <= i + 1'b1;
							CS_Valid_Sig <= 1'b1;
						end
					
					'd2: begin							 
							AD_CSn_r <= 1'b0;
							CS_Valid_Sig <= 1'b0;							
							Cnt2_en <= 1'b1;							 
							i <= i + 1'b1;
						end
						
					'd3: if( Cnt2 == 8'd71 )				//valid CS↓
							begin
								AD_Clk_r <= 1'b0;
								CS_Valid_Sig <= 1'b1;							
								Cnt1_en <= 1'b1;
								Cnt3_en <= 1'b1;								
								i <= i + 1'b1;
							end
						else 	
							begin
								AD_Clk_r <= 1'b0;							 
								i <= i ;
							end
							
					'd4:	if( Cnt3 == 8'd6 )
							begin
								AD_Address_r <= Addr[3];
								i <= i ;
							end
						else if( Cnt1 == 8'd12 )
							begin
								AD_Clk_r <= 1'b1;
								Data_Out_r[9] <= AD_DigData_In;							
								i <= i + 1'b1;
							end	
						else 	
							begin							 
								i <= i ;
							end
							
					'd6:	if( Cnt3 == 8'd6 )
							begin
								AD_Address_r <= Addr[2];
								i <= i ;
							end
						else if( Cnt1 == 8'd12 )
							begin
								AD_Clk_r <= 1'b1;
								Data_Out_r[8] <= AD_DigData_In;							
								i <= i + 1'b1;
							end	
						else 	
							begin							 
								i <= i ;
							end
							
					'd8:	if( Cnt3 == 8'd6 )
							begin
								AD_Address_r <= Addr[1];
								i <= i ;
							end
						else if( Cnt1 == 8'd12 )
							begin
								AD_Clk_r <= 1'b1;
								Data_Out_r[7] <= AD_DigData_In;							
								i <= i + 1'b1;
							end	
						else 	
							begin							 
								i <= i ;
							end
							
					'd10: if( Cnt3 == 8'd6 )
							begin
								AD_Address_r <= Addr[0];
								i <= i ;
							end
						else if( Cnt1 == 8'd12 )
							begin
								AD_Clk_r <= 1'b1;
								Data_Out_r[6] <= AD_DigData_In;							
								i <= i + 1'b1;
							end	
						else 	
							begin							 
								i <= i ;
							end
							
		   		'd12, 'd14, 'd16, 'd18, 'd20, 'd22:
						if( Cnt1 == 8'd12 )
							begin
								AD_Clk_r <= 1'b1;
								Data_Out_r[11 - (i >> 1)] <= AD_DigData_In;			// from Data_Out_r[5] to Data_Out_r[0]					
								i <= i + 1'b1;
							end	
						else 	
							begin							 
								i <= i ;
							end 

					'd5, 'd7, 'd9, 'd11, 'd13, 'd15, 'd17, 'd19, 'd21, 'd23: 
						if( Cnt1 == 8'd12 )
							begin
								AD_Clk_r <= 1'b0;
								i <= i + 1'b1;
							end
						else 	
							begin							 
								i <= i ;
							end
							
					'd24: begin
								AD_CSn_r <= 1'b1;
								Cnt4_en <= 1'b1;
								i <= i + 1'b1;
							end
						 
					'd25: if( Cnt4 == 11'd1049 )			 // " Conversion time "
							begin
								i <= i + 1'b1;
							end
						 else 	
							begin							 
								i <= i ;
							end
							
					'd26: begin
							i <= 'd1;
						 end
						 
				endcase
		end
		
/*******************************************/			
 	assign Data_Out = Data_Out_r; 
	assign AD_CSn = AD_CSn_r;
	assign AD_Clk = AD_Clk_r;
	assign AD_Address = AD_Address_r;


endmodule

						 
	