��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�s8�R�	�}����pn�R��}"6�l�:���;�g؞U���T��ײ2��>���^k�/7�?1�(�c��ߘ�]���<�j�C��`��L&`^����8��U�Z봣��D��L���_�L�3��0I}.�ANMs����C^�cS���N�w	*D���y&�f��+K��[y��ڂS�O��6b\U����/lt�3� P�;��1�-��⫯g*P(�C#<�:z����uP!ߌ��˼�{�&��ѕ���jǎX������n�q5�(�+}c�)�Y¹w����HNx�IL���om�Q*���T�K��͛�����Ŧ�l�N�`�ě/:cї��������qV��6���d�e������2��zEI�Ý�M���A)a��4�D�h�1� ����;�Ӏ�md�L�aV���o�C��ɡgJ����f�P��_�v�h��`O��Ftl/�~8��Ș��<)4�H��vE-,b����Ǘ�Y����<�4�X#�Mwn��A@�r$�ȭ��J�w��<#�+�[�}��|A�Ww�=�d���Fz�!�`�(i3!�`�(i3�<VP�b� ��E����q�B�^��7ص��s�r�X�<\�t7��s���q��cW�sn�;��J8�����3(:�QuK͖!��x�	vy��s^�&���Fz�!�`�(i3!�`�(i3�=��W@y�]�� �OׁΫ3݁_��޲L�&�V�.Ю ��&\VI`,�ʺ�;[��+$�6ﳌl��t�1��꧄�c����E�zy�զ3�0�j,-�q�m��c��!�`�(i3!�`�(i3!�`�(i3 ?[n�:#G٪�t6�yG�?� }[�KO[2vj���B�N� ��b�FP&ׇӭ��!�`�(i3!�`�(i30R��=�El����W\0���JY���y�!��_��0_��hd�Z��N�T?wׇӭ��!�`�(i3!�`�(i3p=�n��ɬc��WN�����<�FxNߡ��IB��<W� g�[�ܰ0|]<w:���G]Fň��h��<�rE��"7HI�S�k�,�B���,���}0xs�Җ,G����Fz�!�`�(i3!�`�(i3tk��mrW^~D�n��������t��p�O%�+�}mIƾ�Nh�m ͠c�|�]���!�`�(i3!�`�(i3H������gf���)�:	<�J��I�s�(�ߜ1�*�Hg>pu�y�jI���뺨���!�`�(i3!�`�(i3�K�Ǔ�\=RJ��z��"��:V������(O#�e*L�E�w�̙	,N�y����~p�7��w��b��rH�>�S�6�0RD��}��b.�Y�PG�(d{��8ѭƦͯ\�Q~!�`�(i3!�`�(i3!�`�(i3L)+l��n�����<�fi
�׋���1�r�63#d�ׇӭ��!�`�(i3!�`�(i3�ݐYs�����'t-/�9D��}��b.�W�BV��(�ߜ1���ccnh?�!�`�(i3!�`�(i3rK.��=(M($FO�X�B�ei���s�61%=��+��>�6AcUgE�ϧ������c�$ׇӭ��!�`�(i3!�`�(i3T�[9�=D֦�ccnh?��sp���(�ߜ1�U`�V�٘��LТ��-������LB�����ɧ���~O�kQoZw�ןLYsȸ�"rR!�`�(i3!�`�(i3]��g��a�5~e��T���c��~$s�c��0ے���(q�� �0���h�)���Y䋇	���1��/z_�����h�[ѽ
�O���6��2�k4|��1+�l��r�����<�>�y&�E��}�y��X2��6Z)!�`�(i3!�`�(i3!�`�(i3ZHm>��.;��L�Oɬc��WN������J�A|������l"9�ۗ��!�`�(i3!�`�(i39�O��F�=,�m��B��sp���(�ߜ1���*ȑs��!��z��A����\�K�y؄@�!�`�(i3!�`�(i3��+�t2���zЊA}.��ccnh?��I,�D�y:#9�]�B�-����;���ԝ�i�Ҕr���7��Pgen�MS��5*��8��i�c�g���H�!�`�(i3!�`�(i3!�`�(i3��o��d<r	�%\*<B)363�8�.D�V�6�˅�ٓ� ˖%*����ֿ����Fz�!�`�(i3!�`�(i3}�E%|0�WJ�Slm�m��}����.HI{?a� ~>>ը܅%Gbغ���:�9��#2c/������=pds~��E&����Bsȸ�"rR!�`�(i3!�`�(i3c��N�wC����P�B�/.w�u�$f���܃n��]ȟ!�� !�`�(i3!�`�(i3!�`�(i3���C�RgҘ�I9�UC�*&�+�eؐ�����!��B���k�c��`�	U����f�7U�i�#!����P�>+�va��2u<�F�x��_���RQ�
�0��,��X!�`�(i3!�`�(i3!�`�(i3L�E��1I�OfUA`���B��ҙ����WH%���ܜ?n昼�2#:� c��(�U��;���-?}`�I��d`ȯ~��.S�M�#0NUD60L�(׌����Ƴ�����4=����f��b�+/ �M�p k
� �,�i!�����"��e����l�5}�
Z$��9�jw���9�ȭ��J�H�M ��,J�l�/�I5@�k{��� )<`w���'挒_�>c�?��ț�?� �عNUD60L��c�6�fSTh��\�ڰ���gLE�z�:
C=�!tC����ı��#d�F�[��m�O�h|���*c�M�B��; ,@�� T���,�� ����]P{�u�$f���SH��{?a� ~>>ը܅%Gb�}$��vk�,�ŭ�O�V2y/�q4T�An�� ���T�BQ���n�n|s�)>ΊՉ���6L�'�1Q��!7s�9��5�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�WOtl����m��c񃰮��^�3�Z>�=�G	�L�UGj��o��]v"5[�Gj��o��Y����6F$90�H1�����\��Hv��3t����k0e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���y�A�T�3Vl�� �̮��I�#<AuA1����v<<,� 2H����QkO|V"��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hͥ<#���vSB��n
HDW�Gj��o�l�����CGj��o��]v"5[�Gj��o�z^Fh&�ȕGj��o�R��(�.cGj��o��(���H�Gj��o�>�N�)-H2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�b#Ӡe��?�F��&k�ZV"���:��#tC������s�Q�_;�"l���c�a����9�ĒTC��0���^S�kC�"�Z<�
�#*t�uADa��?4j��a����2�˴L�t#[����p������*�۽�.�jI`� r��F'�J�|(�����	x]�V������g��Z~Y��]#�]E���4������D��a�,F�7&�����pN�Wu��w)�S���f��^@�~篟|�Q�M�u�c�.C�g�dџ�_�v%��O��J�O�� 0�^"R��#'5��i���~+�lX҉ys��3Tb�����?�����$��w���މ�r�O��C��0��QP路h�����G�/9��g��G��������!�zg�Z�$�����j{X� ���
� �AH��1�����Cn���ʯa9̷�
�Xg���e�JrtΣ|Y���%�����φ��~��➛����T8�{��3!Z�*_#a�/����i���7�`ѡz��9���vo���Q�g����#$^��j8HQ��X�t�q���ѧv;��gf����)F�Z�u6_���͌�<�vd�̪?�d���&��P�>�� ?[n�:#G����8
B�ɹ�`S´ c��(�U����	x]�<��O~��#?���/��di���� J���<���&}Xa���qd��.�wjX5D	1%���n����k�8���҆�|n����﨩R���i&��a��fx���$�U��"�>�q�ax�MU�٣�R�B;����4G�n�?�`7�K�|���g�3] ��Jkŏ��8%C��c�S+d��t4�f%N�XG���\�4�s�q�=Q��xY��݅ 0��|�~���nM�bb5�Sd,�ϱ�ϖe��!I�I�� n "<W55��XR
ئ�v�5ܗu��S&ϊHF>iDj(���ʇ��p��x+65�p����o L�"��\�4�s�q�=Q��x�)�����|�~��wU�����Sd,�ϱ�ϖe��!I�I�� n "<W55��XR
ئ�v�5ܗu��S&ϊHF>iDj(���ʇ��p��x+65�p����o L�"��\�4�s�q�=Q��x
�ԟ�d�F�D�Oo������o?�M��;]�;��
<�����&��*�_��l��f���<zT����H��6Ó�KF�vw�}\yȺ(��m��A� c��(�U����	x]�<���e�0�9�(��`ݓ��� +u��Ipc9�`s�S�͔�Rټ ��߷��\�4�sR���i1�8Y�&�\���p�h�%ģ�l�$9Ř��W(�1���z���D)���pH�P�SyH�O(ٛRF�",�uJEA�����X�(c��k�8���҆�|n���u� �(�eg>��rvp�){�~A �ѕ�����aWfL1�;4�zu%�1<�$z��n��kF-�F敪29k~��e&~�:u��w)�S��X3���7��Mv�9����Dtr/���zbl�џ�_�v%��X�'b�mh}����N�@N�����N���6[�'�&�' �>�u��8�F�D%� ,R�w]�y�ljrHS�w�MH��j���r���+W��YJt�,�y"r� J&g~���c*& z�s�ђ�B�~f��0(�/��$ }2����T���Q���!i��ӯ�02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc/?�s�m/C�Ѽ?��Q2�=W�֯�^��N�&��^˻f��	g�y���}�ZC��aNvA�;�m�\��qi��p�7���I�4��ʆ	��i��p�7��Z鎬����~x���i���;t˩�e�J�4>��1lD�J8���=Udq��D��tw:g+��T��d^��_|��3g�ݜ��s8[Z�`
5��*�z�������D���J7"$�zV���a��Αo��p2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc~����������0��D��L���_�L�3��0I}.�ANMs�����(�l��|A����S��������Ǜ岦�%I^�����зq8�Ј$�F5k0B�����6q����"� _̍�����b9����4�6�t��pf�,�-ެѨ�Qz�����%Ah�%4
>��XP���i-�9c��G���������Q�^�y�zL͊�q��� ����{7$0~'��&\VI`,�����l0��F��jT�����N�i��Ń�b�YL��&\VI`,�n̈́�zL͊�q���$�F�s+���!,�U&��/�,�#�H�1c����O}����g�a!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3f�X0����ߠ�p���R*��7��As?~�F*�Z�"1���,��8�-Zy?X�-r��|ڑ�H���o���&�t.�}�?��E@��j�g��o���7�"��%��^[Ό�������7�ܥ��2������֪zw�&��Rb��Y�W��T�ߑ"��������)	�8V���C~��m���4X%���'�4ɀ�!�`�(i3!�`�(i3!�`�(i3!�`�(i3�� л�7�lcR�+�ye������N}"��5���4<լF<�gH����ܜ?n昼�2#:� ���3�ҺIÙ=�H%v@����f�7>�����D/͘B�N�pS��Y���8�TP���cӄ�=��}2M�; �������@���k��l0��F��jT�����N_�G�*tUL(\Ӧ�H�W�h���Q�#<4^�N�By3��<�]�!����M[��ǢR�����Y%T��BPe.��xu	�>��l%i�-��!|�|~�?�����2��p�c%��C���B��+ Hc��Et��q���U�C#/<���q���V�^��nrm؊(�[��N��>&S�XQ���t	M:HZ鎬�����	�7 �#��$J�L���.��,��]���>����C��(R\֎u���L�u��7G#+��\w��0](@X~�H:6�>u�t�a��(�
t�ژq���U�[��N��h����MԘ]2�y�Z鎬�������(��� E�����(J�f����ߑo�1��� ����P�7� ^�V]��}R�wX���|������kxu�2���HF3U����ޚ��@V�� ά����
L'���Xw�j�7����w�K��ݑ�][HW��W���֨g��U-�e�,���6+�=�B4˖ב����E��@IE�U��*�QN��� ]���f�fx��V$�w�I�?g�f���\X�<����8��UWJ��)y�S*���
���<�s!�Fr忒@2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc	~+��*(��z�jv .
L����1�:�Ω�s8�R�	�}����pn�R��}"6�l�:��\��,�֗q�Z��y���D�I{�����U| �Q�^�y�N��B�)Y}�
�?�?�����&*ì�u"4�JHn��z���i{8�.�@�p+'e�&?~�ő%Ah�%4
>��`���o�)�`E5��1ig!�E����FZ鎬�������(����F�dH�/�R��(�ߜ1�D�P�E6���2����.��c��:KY",oMG~捼�a��%"'���Xw���,D�H�p0���U�)3�B6�n`5�fK�\w��0]b!��u��K�&�a���Z�����]�!����w�Հ�b02�O(�`ʂ粠�+�J���q���U��@����gG�U��5f>U3P�7s�9���o>��l%i�-����]��O�M:R	�G�L3cfi����hD�v�l�Ū�TD���)T&I2WM�vT�V��|�������c�A�L'��~�2�?�B���N�gl��ܬa(􆿳���2����.��DP֞ E2�DZ���ǘ�g��O�M:R	�4>U����������bp���%~����	;��Hlό���.�	����$�qcW�(u�" Oag��đ�O�v�(R\֎u��O`ALS��(R\֎u�z8��oSx|Nb��'1-Y;�e�O�!�ўC�k����}o�`�������i��.����.��$|�;�Ojz�>��.[[|�;�Ojz��o��3�|Nb��'1-���9�~�p�@V�� �<z7n-��8�8�rS�Z;#��Hۭ�#✲�@�ZF���X��ߊ�ֲ���ܜ?n昼�2#:�g��U-�e���H�V�R���Bk�d�#✲�@�v/fu����1��� �U��֜��3,0=]^	�&���忑������Ho��'�\�n��F����Y:�HCaIMl��ù:�h�aT��3G?�d���&�8�w5+�uh����M���Q>�����T��_
fg��* ��>�:�;�Ղ��"�[(��K�I� ���	�Z�kfcv�q21�ю�=2�L-�$��^)B�!�`�(i3�E����Fxy0�u��?�;���]�Y���v�岦�%I^:��%9&���;���EWrr{�"���!�`�(i3,ԯ���gnņ��#�b��~�26��\��Y6�ޤ�p2�]����+�J��Y�{'%s=ͱu���˝Sz��E�4.@�7��y%%��`y���ֱ�q�����2�w�]'�-Q?9�!�`�(i3���#] ��2N��n��k�@7���K�)�Z3"�,�>E��ʆ�In��t��+x�r����l�©�oo�@L=��\�ߜ7�ܥ��2�����r��%u*w�A�2N��n��z6��@�
�zS��jj$����c���+�J��YV5����4���܂��+x�r�w�c*��R��E���!�`�(i32c<���z�wnB�K���X��b ��b�FP&
�E�6�g�!�`�(i3*�,�3��FP�?��{	%v@����f ��b�FP&2���p�!�`�(i3*�,�3��FP�?��{	*.�PS��� ��b�FP&��$"'�ь%�"�Z1��X��ZG>��|��4Q� ~��d=��¾ȼ\���F�`y������T�8k��.ͥ�H�RtV�^	��K,����z�щ�%H�&��h�d`̮�ӋH�RtV�^`��M��v�Gꉼ7��b+}y[�y��j��k6Z�٬�[���e둼�;��,۽���ݚ�Н�V	��V}>�O���(Cq_c�!
�T�r�5�.��J�޺��:p~	5@�=���
�!@<Yɞ* Ϗ�������l�������"�,%�R�H�Mp�Gt����*�.U怺�ݚ�Н�����a�~9��tf��!���z�щԑP�מ��!�`�(i3�q�	��c�O6�k�v�"E&��� �=+ӓ��#!�`�(i3~�`cC�4�. 9ݹ���2esdo���}Dq�f��r'Z1p8u̀A�p���gRI/�|9��zD�	��x��ݚ�Н� �ԣ�e���P"���=���gRI/ӝ�9��,��5����Иy��j��k~᭜�aG�vSB��+�E4u{4��ڳ�&:��b�}�D�ɸܢ�hJV6��c�O��͜N\�𱍞3ƥ��kE�r X��}Dq�f��wbk�$���Ѧ��*n��뾦�!�`�(i3�<�W�7k��#��}Dq�f�R�͢��n-���!�v�i�9&� 2����}����e�]�Q%�1FXM升��	��m��{ֱ@��ݚ�Н�T�zS>�jA��x)�%��U.V�ݚ�Н�T�zS>�5�xo.`�z��̗��岦�%I^<�5
���d#����*�
�:qEp�;�P�t�5fĉ>99��A0ok��EOJ�uxm�Q�Q,4�x����E2b�z'hۉ)K7͍���E@�����}Dq�f�����0��Gd�~{��)P<�ܓ�Y�99��%8!�`�(i3��ic)�̩ƍ2���l�����g�Z��3��a���!@�f")u��r��$XR�QܛOcOZail������&G����l���}����O}
��g�-����� OLfq�n7��
�����VPYu��r��a�}�$�ϔjZK��#��_�?�tT�_�X�p�c�ݚ�Н�y8�:����G� �X>���\4T۪�؉_�'���~� ��S6��ح�	��7ص��s�k��vy�e����O%���ݚ�Н��]���`T�fD��j���eK�	�$V�#o�]�ʄ�;4�zu%��XW�G�<��g!4�s��(R\֎u�eK�	�$Vͯ���VPYu��r��!�`�(i3��֖+�){?a� ~>>ը܅%GbNÌ�Y,�u��r��!�`�(i35�����}Yms��/�u���4���O�>�k}�r�,0=]^	�&��|�B�����Yk��!�`�(i3�wbk�$T��8$2OU�1Q�\��^����!�`�(i3!�`�(i3���vO=�)�`t�`v������}� h�ҩ�!�`�(i3���y��lD��&	;sзZ��F�$i|�D�yX�ݚ�Н�!�`�(i3���iL�z�
�X�nZ��3��%��|�)�[TD!�`�(i3!�`�(i3q�\E��0N�]|-��{��p��N�m�[�N��}Dq�f�!�`�(i3�	��x��ݚ�Н�!�`�(i3����a�~9��tf��!.G�9^&���}Dq�f�!�`�(i3q�\E��0N�]|-������:Y�{'%sk����w�;{�'8{1�'e���K��!8�#.��#��Q^�MY:fbmDF�!�`�(i3!�`�(i3��Ě�����}Dq�f�!�`�(i3;�E����hQ�N���QK2�(T4�~$����-^A�{���}��n�����o� ��@H�ٗ�'Z!�`�(i3!�`�(i3�{���e�������r����Ϟ�
��-��HF!�`�(i3!�`�(i3��Ŷ�O����Ѧ��*������� h�ҩ�!�`�(i39��n�7�Y���X�q����;q���Y�l,`i.����!�`�(i3!�`�(i3���F��O��ݚ�Н�!�`�(i3�?�JY�)�Y`��jD4�ݚ�Н�
�:qEp'{w#/ B!�`�(i3�wbk�$T��8$2OU�1Q�\��^����!�`�(i3!�`�(i3�R'cf��i�X!�!D��(J�f�x��2�+�T�\ ��[��(��!�`�(i3!�`�(i3�w%˕1�,��"<���t X��ݚ�Н�!�`�(i3�� л�T�â�v�+�X��^r���C)T�!�`�(i3!�`�(i3�y�MP�<�����$��㇟�})�1C���.j�!�`�(i3!�`�(i3w�����A��ߎ�x��y�2р�����T�Qpr!�`�(i3!�`�(i3�����!�`�(i3!�`�(i3�]��/ݐ���n�@���^����!�`�(i3!�`�(i3w�����A��ߎ�x��y&k@C�Ɨ0z�cULE��K3�j����,�9��tf��!�7>�����ǚr��yݲ�Z��*�!�`�(i3!�`�(i3�5ߧE4��!�`�(i3!�`�(i3�^ ،�X, ؖz���d9=���u��r��!�`�(i3!�`�(i3���gRI/J�a$�Y JP�l��"\�$���!�`�(i3!�`�(i3��Ě�����}Dq�f�!�`�(i3�?�JY�)�Y`��jD4�ݚ�Н�
�:qEp�;�P�t�5!�`�(i3ݑ���&�d>&S�XQ�<F�ڴd�?D�8��!�`�(i3�5ߧE4��!�`�(i3�����!�`�(i3u�RV��,)kJ#��t��$VĶ�A�2n!�`�(i3��#�a�Ą��$J�L߉����<<��lp",oMG~�>y�pA��M?��y�!�`�(i3��l�^!",oMG~�@�S?�PmƊ��NM���!�`�(i3EOJ�uxm�Q�Q,4낆MC@���1����?����}Dq�f�՝� s�#���k$ !�`�(i3�(R\֎u�eK�	�$V�%��v��!�`�(i3�2��}��E2�DZ�⦫/���bxK7͍��wAA�Ɓ=<�W�.�P�H,0pMp!!�`�(i3���F��O��ݚ�Н�$f��_Ub�F�S�1 ���w�w:�!�`�(i3��Qѳ$G����C|
�ݚ�Н��c5ew���$J�L�l:�
d��<<��lp",oMG~�>y�pA���Q�Tq|�;�Ojz�$�AՁ�';��#j�ݚ�Н��99��%8!�`�(i3��ic)�̩�?D�8��!�`�(i3����0��Gd�~{��)P<�ܓ�Y!�`�(i3EOJ�uxm�Q�Q,4�x����E2b�z'hۉ)K7͍���E@�����}Dq�f�HN��R��bP�63Z�tHN��R��bP�63Z�t��Ě����E�i�m}6O�D mWN��ܐ�}��y������h�G��2�IZ��O��<�� ���`�ϦE�6����ѹ��6[gb�r	�BS�eL׸�n��&v�M�,!hޖ�A$�P��O�@יߌ��omq�:Fa�7������A�ս��*��Ͷ�2��i�U���e��d9=���u��r����z��A�����**,n��;c���k+Q�h'�Ȝx�5W ��̫(� h�ҩ�:
��x�{�\��N�Ś�-����;�jmT�#�(R\֎u�eK�	�$V�#o�]�ʄ�;4�zu%��XW�G�<a��o���H�RtV�^��#�a�Ą���*�����:�I���Oj�\Ʊ�������=aS�H��ݚ�Н�џ�3~�l"+�B-�D^օ?D^��!�`�(i31���~!�`�(i3?�����&*�K��d�N$���*���b��~$�!�`�(i3���F��O��ݚ�Н����F��O��;b�-�2��;�P�t�5$f��_Ub���uQL+��φ��<�6�?�����&*Nۂ�k���V��QK��5e�Il�,����~��}�m���ޙ��� b�	��6��*��1�u��.t�5�M�1�>�0�؆�ʷ����{d�T�d�U��o��_�Rv�䩲$����#��i黃tx�Xg��(y9��^$�xKw�66l8���x�;���EWrr{�"����a�\�����fZ���o ��b�FP&p�]f�"v��os�z���+x�r�s�*�I�qcCl���<�[fc��RC����Z����1�����:$�:��q� ��b�FP&��N�T?wg_�����A( ����_ֲ��mŹ����q��iI9�o«IX0F�M��(G0����2C`����"sS<GYqcHTX�';��#j�@��v{�G�n�c��	nK� |�>��� л����!ɿS�Ĕ�Z�_d=
&�|p���s�-k�9��V�9����m?�Q�����z1h�'��H��/��@�ذz���:B�a2�dZ#'��� h�ҩ�T�zS>�����i֘JmՑ�hS�nJb�G �<��hCZ�� �0����pX���.I��Ͼ��\�qj&�G�;�jmT�#�&5�/h/�[�a��O��_��-����!�`�(i3f퀔����W����Qy +߂X}����e�V�~5�f�j�s�B�4�x��w���0v
��[H~����}Dq�f������!�`�(i3�����i�FQ+��1%��[	J��;��}Dq�f���Ě�����}Dq�f��5ߧE4��߆�p�h��d��JXl'�T��~��Uг�|<;�jmT�#��"����G��Hb� h�ҩ�i|�rBY�",oMG~�>y�pA��x��w�����$J�L�l:�
d�^��.�m.�
�ɺ%�K��^/p�O�޿M����eo>��J�M����!�`�(i38��A�8N�;���n�c��	n�T�TN��!�`�(i3����m?�Q�����z1h�'��H���b=�W!�`�(i3�@J`�]���xv�����C.�u�X��I�ՠ���Kf����<��ޠn!�`�(i3a3@��[/�L��O��pE�<l��uE9�+��!�`�(i3{[�ב�C���#�'4v~9��c�	?�N����!�`�(i3�5ߧE4��!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN��Ě���aT��3G�IX0F�M��(G0��:��1��F��A���9��d��z��w��G�$U����KmU��@B����,\ަ�It��bF��ԣ�����E2"�+��O�V2y/�	p��+M��ѹ��6[��{ֱ@�gp��{k�M�Ax]�ǒ�x�aRom9�����*�/l������;M£>�2���w�c*��R��E���X2zӼ<�z7�g�+���ֹ�͈����$�Qu��`2|`Kr�|�KT�Y��]��$�]�#A���+x�r�s�*�I�W2��H9��d�������|���{�����~�26��\��7�8�7^XX�<f�K��\�v���+x�r�u�#��nt��F�z�8# ���3�Һ��7U��s���+�^n=\f�5>���D�����d��JXl'�T��~��Uг�|<;�jmT�#B;i�L�jrq�A��Дd�8��k�S��?�9�7#1=��*�����z��](g����>&S�XQ�u�j�fKç<<��lp��N�DNlvr5�Dѯ�p�\ì���uxrBZ@2� H���YCթ��8>&S�XQ�������;Ȼs��VA�ڦ�c4�L2A���b�YL��&\VI`,T��8J��6��˂v��la1�ݚ�Н��� л��5����`K ?[n�:#G6�aI�[��!�`�(i3��N�T?wX����0<�Y�{'%sk����w�;F}���V6�����a�(�ߜ1�3�N���[��}A?���`ޘr��!�`�(i3)�{6�U��ʁ���MյG
~�	>�3��Y$����y��lD���g�{�� ?[n�:#Gb����HA!�`�(i3�Hx&6��ѥh���>�
�E�6�g�Z~~���<�:5A��p�/��@��R��E���4T�Sq��{����[��d~(N�����o������P];�!�`�(i3�;�	��o�2P`:vS��h̥�5�8}�gB~�RǏ˨�g��H�����?�@,��V�'vX[������?1�lm![����{_a\F!�`�(i3�GI�\�0�c��v��tz���*�m2ٲF���ؑ�c�ݚ�Н��� л����ؑ}2O�V2y/��As��s1���]/���^��9��m��H����+��l�t�==�SD����r����<�6�Q=�v��6
R�>���:EW{��.�8�ݚ�Н��H����}���yb��Ҁoŧ�˺�&\VI`,9��9dJ�!�`�(i3Z��JP���K���&�G�T��}��T�#_�B�ݚ�Н�fĉ>99��A0ok��!�`�(i3�ج�B��l[�Ƶ��p�����Ѧ��*G��Hb� h�ҩ�!�`�(i39�F ��T���$��w�kK�o��oW{TT���.��k ��!�`�(i3���lS���|�+^/�����������p"3?K�[!�`�(i3}��Z&�G��bDe��Z�9N�^p"3?K�[!�`�(i3;�jmT�#Qi�d��4�T��ј|� h�ҩ�!�`�(i3 �ԣ�e�	P��o%z$���5gK!�`�(i3;�jmT�#�R���"'��h芼�o�ܺ���N���!�`�(i3!�`�(i3��yl�6��PiA��t���y�c�(�ߜ1���-����!�`�(i3!�`�(i3�����i�I�p�dQ�I��F�z�8#[�Q0�M�!�`�(i3���%>�rGO�D mWN!�`�(i3���%>�rGO�D mWN!�`�(i3HN��R��bP�63Z�t!�`�(i3�����i�m����pe�'���Xw�j�7�����P�|T�O�޿M��}
Ĭ��S��1ig!�l�-��;�:5A��p
�:qEpMH�%��LX}��nM"��N�T?wl��a�.����J�4�,��M�9]��-����!�`�(i3U����ޚ�^�OG(�((�]�!��	Ǹ�y85��8��,	i� ��V���;�I1��N�T?w���[�����qE�N!�`�(i3�� �?Ct(����ۘ�%��v�V��Tk�w���g�{����7C.9�����b��n���S�P��~�]��%E�!�`�(i3��w�w:�!�`�(i3=�'*��{+�d�C�U=�ZP���m"Wm��|ɟ)�����I�!�`�(i3�����i��i�+�؝7�q����	Dai�4�d�C�U=��[�[@�B!�`�(i3U����ޚ�y�e`��&k@C�Ɨ0z�cULE��K3�jAԢ�a\�%o�P��(�cR "�=���y�pkv|p!�`�(i3�y��j��kb��4��;J�[��?�8=�V����Vp�ܬ���������Z!�� j�5�p�mҷ}["��4�}���yb��uE9�+��!�`�(i3�5ߧE4���ݚ�Н��� л��g��1�Eղ��>e<�6�Q=�$�lӪr�gf����7� �9��|�_6i���6��V(pyL0D?yz��������[jHN��R���
�Ŏ��HN��R��bP�63Z�tppE�"f�;�P�t�5��/z*q+߸��S�Ȍ���=g�6� qM�[���6<���ὕ?�5�e���Jm�Wb�#���)��}\yȺ(��m��AՄ~����p�����%����:��~D(�kw���'���WŌ���������:n�3��A@�r$��,�c�S�s��ǿL��D�ݓ#_}Cd�_���S�# [�T6;��|B��� OD/=3\H��8~e�o1n�K�S>��zL͊�q��sM
������S&ϊ۩<�r�[@}	�׫�i3U��P3z}�&�dLG���6�C|�����!�wc����M��7��o�Ǻ�j����2���,�ۺ�j����26����$K:E��]��8�]k�Z_��ݷ�pB�aZ
��=��ݷ�pB�a�e�����0��èV�S�D�m̲9��4�φ��<�6�������y�:Fa�7��Ɨy�"c�Յ��og�ѓ�+g��U�Q��$�pٳ���T�B���ќ�}Dq�f��N��[r���X��ټu��.t�5�M�1�>�\�l0�?<�v%_��,e����Y��˃#�c@X��Q���_�A�����L2���gRI/}@�̵0z���-8p~�����O���}���Ȓ�/���
.�/��H��m[��k�(+;���%�4��%�p�!o�{^��w��b���u;�`@t�{f�U<I�j��ޓ4�Y�qHJ��ՒǸ'o��j��ޓ4�}Y<� �х���W�w	4V��߼��:�JKoW��sj�וN��j�K��R���;kUZtץ���:Z{G�id'�t��]��N\�Sdb��)�E3	��D!,�$�5���y���r	�%\*���l�l`�x��c��bƑ�����߆�-M����k<�6�Q=__�n3	r�-�@�3�m�j8�0���R|�
K&2��m�qH��G~�U�Q��$�f�Ç{˙+�B-�D(���27:����Kf��w�n9�gg�;�?[��t",oMG~�>y�pA��x��w�����$J�L�l:�
d��o�������3��a���� 3bH2ȓM�Me��HcnD��Z
�7$���ɟ����x-�	B(�	<��	gvӯ5 � � p{%AN__�n3	r�&���"P �h7DP"G�wk���U.+"b4��ϗ�](g����>&S�XQ�u�j�fKç<<��lp��N�DNlvr5�Dѯ�/xR��\&4��Ȝxڸ�c�K'�<�6�Q=Z�'�!��h�E���bK���Ų���R��-�	B(�	<��	gv����VGҺ�J����+�Ü p{%AN__�n3	r�&���"P �h7DP"G�wk���U.+"b4��ϗ�](g����>&S�XQ�u�j�fKç<<��lp��N�DNlvr5�Dѯ�/xR��\&4��Ȝxڸ�c�K'�<�6�Q=Z�'�!%<�e�r~bK���Ų���R��-�	B(�	<��	gv����VGҺ�J����+�Ü p{%AN__�n3	r�&���"P �h7DP"G�wk���U.+"b4��ϗ�](g����>&S�XQ�u�j�fKç<<��lp��N�DNlvr5�Dѯ�/xR��\&4��Ȝx�����\�JW?�;��Ɨy�"c�Յ��og��p�n��n�ɈDf%��U��)������|
l ���RK�*��gB���~���v)�ww��Y���d�G}%����3f�15mo�����Yk���K�&�a�W�^�|��/��kOT(@X~�H:U�)3�B6%��v�ڪ!�x=�FZq�%��\�m��d{��A��(*�O�q��
�/fղ��>e�p�c)C�+�B-�D(���27:����Kf��w�n9�gg���-/a8!�`�(i3�(R\֎u�k�n�=��"��ӌ�r���%>�rG�@�	������6������X��.T��;�jmT�#?�����&*��,Յ�1tSjv���+�t2������gZ�_v(���?D�8��HN��R��F F�E̠ʁ���Mյ�#���6����$K&U�)j�S��#�a�Ą���*�����.��y�� h�ҩ�ݑ���&�d��b��MF�̃��H��}Dq�f���Ě�����}Dq�f��p�c)C�+�B-�D(���27:����Kf��w�n9�gg�8�fk!�`�(i3�(R\֎u�k�n�=��"��ӌ�r���%>�rG�@�	������6���(�wJ<$&o���՚�jT��;�jmT�#?�����&*rB�WD�{͘6��q����1ig!��'�W?�����&*��,Յ�1tSjv���+�t2������gZ�_v(���?D�8��HN��R��bP�63Z�t��#�a�Ą���*�����:�I���Oj�\Ʊ�������=aS�H��ݚ�Н�(@X~�H:U�)3�B6n��뾦�!�`�(i3�5ߧE4���ݚ�Н���O�������ϒ!�`�(i3�K�&�a�W�^�|��/��kOTݑ���&�d�+��\������{���}Dq�f�)�{6�U��AL(�z��?\�z?Xk�$�)�vx	��$a�O�<F� ����t�td���5��;_��8W�w��fDy�mH�6�\kB�,F#K`'�#�v�*���{�y'��BSBw�>�(�s�=e	6'���3�!SC���"��y	��Mn{�8�
K��M�8Dp�_xغ�#��@����+��O�r!�J��:�����(R\֎u����>^17ӻM�{�|Lɲ_TGt�/�����>w��jVѭ@!�`�(i3!�`�(i3V[B�5�m(@X~�H:U�)3�B6��x�����Xz�Yx�P �h7DP"G�wk���U.+"b4��ϗ���jVѭ@!�`�(i3!�`�(i3V[B�5�mw�R���y>��yС�M��7�-V�6��1myt@w�	��1�eq�z2� �X��Ƀ�+$&�F�6*g^hI��X���(EK�3}<r��m�U��l�@E���af�P
WF�j���φ��<�6�@a� ����C�'�ąd=��¾ȼ\���F�`y������T�8k��.ͥ�H�RtV�^�	�%1A�"��ӌ�r�k��^�1��dc�@c�����h��-������#�a�Ą|�;�Ojz�$�AՁ_�mS8<�n�ݚ�Н���Q7lY��)P<�ܓ�Yfĉ>99��A0ok�����F��O�\E�W��4b����A�ձ^�Qb�Up�C�
���G>,Z3���ڥ����Ⱦ-���H�� �7~�	 �b~*��s��(R\֎u��Gj7�uz�Va�irɟ)��<�B_�2���o�����	.4�0
���gRI/��F�3h��V����Z5�p��ާ�����ݚ�Н�{�d"���Uo�A���8�ܩ�ò�CFy��Q�F*�L��!�`�(i3��7I��ك�8ZѴ`����ǆ| c�]hgi�K�%@2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���j
�D