��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�.�&ʺr����$lw��ܴ"8;�]��;�Iώx�t���E�L#uc��WŬ�+�-ޗ(huUPc�k�u�}�|Ѽ�r�ν��e��eG�I�?g�f�SL�<.w[!�� Q鹯e)�Op$C^�cS���N�w	*D���y&�f��+K��[y��ڂS�O��6b\U����/lt�3� P�;��1�-��⫯g*P(�C#<�:z����uP!ߌ��˼�{�&��lV��n��oNaW��4J�Ś��
��H,7f�t�뾌��ߞ�:��L���om�Q*���T�K����Z�e�g�]��s/$W�o?=4��{0��d#m�sj�]:#���c���`�G�YAds£����&����S�BgV�g�0���ή��M�5���Cd�
��S��6��H4�
� �AH�}��� �Ȱ��-+�T�8�hF�_!�>>��S�O1����h��]3�;���[=�%�
�R�+�hV�;/=�n;i���2_�q�JX�����@�>��+R���RL�a)=�y�~ ���������ߤ����Q�=�>�v�ֹY���8＀�L��q�Jp� ��g������a6���r<����}�a
��{0��d#��翑��HF��eUٻo���mi��*	�ť�.^�i��' 1wH�x�xs��3�<A����2�P`��������~�+��,/,����W >g1�]l�&Y��F}갨y�����# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��`y��f2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�}�Z���ik2)�
}wʭU&H�1��8�h7H�u�ÍeRuw�C?3d,f$�7Q0�"<�F�ٴB�I�SbW�{b�2"���Bpш�#w��s8[Z�xZq��t�1�:�Ω�`<4}��o�r� ��J��ݪ�nX�#fZC��	g�y�+��T��C�NJ���1�:�Ω�A��>s>;܆L(,�TfI�k��S�����ˉ�1�:�Ω�.�&ʺr����$lw��ܴ"8;��M:��;6aJVlO/����\{F˯�+)��ʺ�;[��\�v�W����ĮfA��x�%�ܐ�ʟ�]�AZ��:I�"_��V����p{���,�#������s�0F�2�^���=���8��/��m�����W���9�GW���!��������F�┠�Gj���X��XM��d:p{�imlK:�� +@���0X�K�9D���o�j�0�J�vt�OF��������g2Uo�H�0�{�?Nt�!�ei�P�?��'&�s��Ia�|���+,�)��R�ᑧv0-�(4��AYp/ܷ�Kj�.�J�����;*OZ3$�" ���;%x�6��y�g<.���3Q[����c8?-+eN7��c��;��\�v�;)'gf{H���o)�]rH����8��,�S����'n�^0o��~+�ݗ	��(l��U����z~��;ε��IÙ=�H�S��M�����0)]��w�b^X�P���ma������	�5�V��On+0�l�R<�q��f�}��?��[���-��%Mό���.��_F�k-�v�ј�"��Z鎬����F�71�B��O1��m<e.��xu	�>��l%i�-���6���p<��:�ҋX����>��l%i�-�[b�0<��c��Et�Y�{'%s��.|Z���I7��-5��6��	���`y����ꢤ�Og�ś� ����]�!��	Ǹ�y85��L�@��f�U����z~��6��	�\�HP@�a%=dϖ�i�@O�x�7�hWw�d�pP~��)%�����D��2E�����q�P ڨ��S���Qߵs<��7�m��+F��8�ĭ��{0��d#܆L(,�Tfc1�-���ml�O�� �0w�m�ڍI� ��j'�}��^u�މ\��K��]{���Ψ��F[�σ8��E�ߥq���P��ʬ1H���ih}N�}h?��].�Ч���S1$� �!%��b���á2�7�?��i,��&lG#;�:E��$vi�N;=��c8?-+eN��zʛʑS��_���!+}$|~ïSup�xg쬉� }�����v�WM�v�1a|JHn��z���P��(�鏄��m�q�»Ą �N��B�)Y N��r*�1W�V�bS�-�=q�:�G�c/*��t�	��{��E}��kA���g�AmY�f�aV6�$p��9:6�5F�&� Nm�Y7 �.�AmY�f�e�Tpv�t�	��{����f��r/��5Տ�E`���k.�C��(�d^�ϓ��ִ,w!~�{�xj��V�������j�@�
��_�˜` uqIUe�n
V~$��;*��I(U���v�:���2c���]��	W�����@����PǨ�o*� AmY�f�ʼS]ò
�A��v���%���nJ���}����f�y�6�,���s�M�Sc�j H�1�t�U�:���2c��O�S]^N���U,D�e%�pV���ޙe�����?Zkܼ����Ҳ�(����E�ߥq�X��WG ���v��syu�x�BU�����T�7<�[b%Ɨ����#���Y7 �.�AmY�f��9=�E�n��,��/���
��_�˜` uqIUe�n
V~$�v��syu�铣\Ŝ�zR���b��˓#���o�u�Q�.�c�&��h�X~��6�='����R��zR���bT��l�rG�0�����&[�x�R�"��u���"6���F��O����Z���׏�����Mc¦�.��	���PJ��K�6}�8&x��ߜ��}��c�ҩƮ���開�E��kUȔ�Ƃ�=89����gۮBez����AmY�f�4 T���&�]�F����M��_(����@EM L����`E(�����.{2Y��֗F��^[_�e��IÙ=�H�xI�2^)b��@ŋ��5k.'C���Y�V������p�0ty�P���Պ���pOz������v�WM�v�1a|JHn��z���P��(�鏄��m�q�»Ą �EM L���̟sE<y�t���6���`y���=k�Rm��̬��[�]��z���;�Aė�];�'\{ف(�7���n��T��%-|����A�{G��	�S����p?�z�+��p*���Ŕ���GB�R���>_���[G�_�3��`���c8?-+eN���	;���U,D�e%�pV���ޙe���5ߧE4��(�V�ܼ��������0u�\k|#�>��� 4\j�3������s�أͽgF"?Z�M����o���wu6�Z����Ofۢ��%P7j�7'c�?�JY�)�*vX¸`��ć+叔�$��*'ΕL�tD:��@-�;S5b	B���ddaWL�@��W��]���y�"�V��q&=�a�7�����gP��U��%:��Q���n��j�S����3k��g1��&.��8ݾ+��f�p���#���F�]:���O����	�c8?-+eN��#�"���|1Cv�Ts��E=�����-��wg�V'���$��"�t�
�W��]���y�"�V��q&=�a�7�����gP��U��%:Y�*4<΢�n��j�S����3k��g1��&.��8ݽE�c�t�W.�c�&��h�X~��6�='����R����\���o����"�ϴB�ܪ?EB�>�!��<������GEV�X�d^�ϓ��23�Vw��šB)�Z����-�a�,AmY�f�Ƙ�r��5ߧE4���]��	W���/�zU�=�����?H�
����Ѓ�I 1��6�Ӭ�&�L������)�x��.��p�4�K,sp�#��"Z1�Sc�j H��2$%-���t��B�F�w��$�D-�;S5b	Z=������WE�|������'��ϩ��z4�g�d0פ���H(���Yy7uojr쇤�oZ�x�;��c���X����<�ޚ�U��%::�����=~^5�C���U��%:���3�}@d��=�~����Id��v��syu�$�3\�\�T%��s�`>]ʄqL$&[�x�R�"|�����-����3�}@,��5�S��5��V;T_J��������Lj�����3'��1�P�	�%Ѣ��-m%�u��XJ6��cIH$X�(�J4U%��/�C�_S�䡢�d�N�-ݵ���ď�f5an0	 
�Za`����� T�rg���%�P���jd�^Ι�x���晈�?y���,�Pd0�[X�b\g�`����Wf�חο��Ռ�Ѿ��/@�[`�A��dgbi`f�H���\)�^�!��l�;e��iAl션[�������C Ln��S�W�.�p�2�zgf�z�;qǙ�d��hwMfA�t����bǆhr��(�c8?-+eN)p�D�C|�Q��uMU����z~I-�����)�m��'A>V���"�V-�B��cȬߝ��v�f��'Ƃ�n��\�v�G�y�G� �Ac�N�A���1#%�"Z�n��[���Åޟ6eF���:&x/����Ld��gƒ
�cc�V�AmY�f�A�j%��f�/؞�{����֗F�~;��Yv��\�v�n��l������}�v���Lj��ݒ�Z����r��(�c8?-+eN�I��p�"�/؞�{��WR�`\�n�9$[{^>: 8���@EM L���=�����[<���,Y#A�g��U-�e�/CَA�2
�]��x�}Å�S�jI@�+�{�
�cc�V�AmY�f�^W��.P5/�H��N���IQנF���ϖ�|����=%+]Bo�A;h�F�sZ��;ӹ*"v%)��Qcm h�]�!��	Ǹ�y85�-�)�{���W��_�ړ8���/��Î+,�C[w�4��<բ�]Z�C�;�n8E
;�GI$��ǂcY�~遟k��P���˳͠m�xW��9u$d9�cx�S�����S8�*��G�{ �D���J��8���/��Î+,�C(�X)��t$I+�V�6IWJE�r���秹�3I^�v�[�9q�Y�{'%s�rOw����A�T�g�v���>�֔�=���Jt���wY�$�q
$�үe������hM��1o�l�P��~l|����N���IQנF���ϸ�U��?���D|	�õ��Mn�;��c���XyR�b!����`y���pzl��a�;Tti�� iJa��������ܖAA/���G�c~C�|��m=�L|Dt �PW��a��K�TR"K�g��U-�e(��w��x�ȳ�5�(�T�\ ���|.�TӏR}���tE�U>�f&��'!msR�����׺;˦K��b�Jhf�|�Y$�h�ya�����aU�`�K-����16X{�"��}�u4��d�bR�wX����K�Q�1�R��j}�C���&��vt�3\�ݢ��T!�T�T^��\�z��cSS�b�(Q6D������������C �Q��Y����Qs����[�=�5x�=�C��Y���¡Ȇ%{�;�������aU�`�K-��`y���pzl��a�+��%�k<�̓q�i&.`�]`�?���� ����C �Q��Y����Qs����[�=�5x����E��-���¡Ȇ%{�;�������aU�`�K-��`y���pzl��a��+?B�OA�4�˕gAy.`�]`�?���� ����C �Q��Y����Qs����� Ei�lmZ���98[ƜU}p�<�_�Z鎬�������(������aU�`�K-��`y���pzl��a�8�|P�nkY?`����n`5�fK��0z�cUL��W?vxb���C �r����������ݓ��E��he�C�H)�{� �"�d�٣��c�A�L'�b�F����Wá.��a(􆿳�f����DB�ȓ�iӚ/�N^�������r��1�Z���=� ��j�L�R�^Ƒ���<�3[�Wd�%l1=h��2��+3�n��5�z.�&k�N$
Ҝsݳ+R�G��?��kT֙*��Ɲ���q��/c�z�5T�ۋ����:�NC��qU�PӅόKK�ϙ#]��I 1��6h}�L00:d��;%�u��T�!EY= ��
�����;M������5d�N���
(��sܴ�W��K�r$ɓǃl[�Ƶ�n
V~$����YL���d�gGo��@��]�W�m�4���܂E�g�������(ӈ��Z��&61�8�|P�nk�Bzo���h}�L00:C?�Q䨈硙�t�\K7͍��|��W&":܎#�o�h�d��JXl'�T��~��?u��C@�q2'��8�Yu��"Όd)���*vzwιx� �Q7���$=Q7l��C �Q��Y��nd�,�&��y�7/��i8i�+o{�"��}t��tw�8���/���;�	E�he�C�H���0���G\�=KH�g��U-�e��`��G�9/K��_�&����aU˙����Wѫ���Uh1�:�j,7�H1׏�����M/X*F���&�2Ƣ�IX0F�M�Ks&�eV��	��y���˷�!R�.��>=¡��Lא���!�d���ڹx� �Q7��GL�M���6�N1�J^ ��.`�t�q�&{^n���pN28�QY>��g²P(��>_��f��`;A�@�۰V��`-�.�l��rq�B�3Y[�z��/� ���P"G�wk���91�	m�"��j���U䞃�
��=���b>��xc�1���"��y�X`��_/���	�n��`�D���R:F���Q����"O����n��T��<���,Y#A;��|B��K�l}G�`6\IO߀\{ف(�7���n��T��<���,Y#A;��|Bj��!(�#��B)c�"ü�`0�/�#g�k���pAS��4V}-�п� W��$0���>���ˤ3��g��/���k��Q�D����t��y��8���/�v{��lw	���T8�}���p+��i�~͜b
BqBé��U��֜��3���HK�A��n� _J�/Td@��c�����M�~��~@�H@'X35Y��Ap��E&���?�d���&���Gh�d��؀ǏU�e��FR���'S/�_wπ>jzT�;D���,e"75�E��W��_�ړ8���/���y��BQ@�U>�f&��'!msR�����׽��9\�	Z���/:���lC��U�T�\ �ͭNjX�U�6j�"HsT����'�۪	�}a?�d���&�{Y,�s ���!Όg&W�w��fD���V����'G�+R��K�I� ���	�Z�kfc�0�	���{�c�	�j�-��������I(͂X��WG ��oH��65���D5�|��7�OT�,���p+���������Fb������AYЭ2�2���X0SȗYo.���Pg�,ǐ��؈a����q
$�үe������hM��1o�l�P�u�)�'�m�b�vA`vK7͍��|��W&":#k�˟ܒ�P��f������̀mfF�5.]���^�����p�@��F�KD�Vr[/}>5��0jJ�_/�+�d=i��_��8��GMX��WG ��5��{�3�H��<�C=��~���cO7}�»ԯ�J'>cI��@%B��qĖ7v��\���D��P�)���i���,��V�.o)q
$�үe������hM��1o�l�P�u�)�'�m�b�vA`vq
$�үe������hM��1o�l�P��~R��b��N*�95��{b��vW'��}�D�Tu�^?�&^��9�׍�����u���?�)����^�{"}W;��ܐ�}ħ@�BY���H'>$����,^�_�Sx��E|����_L�f��bkzڱA�e!�.)������0gڊ�e�Ө��'�h�������;���EWr �X��E=rD�f�,��^�:����U��֜��3�T�\ ��������\���.@�w��o2�Y���hu�"=����m��'A>�g��U-�e!ľ2��H��kX��z�*�O8�ZoݮC^eG=���j+�����svy�:������u�%#䦄!L��9�o��!�d ���g����VrAԢ�a\�u��8�qmO;��%YMYo.����-��U��{H�3)-~sEz���O�cSS�b� �C� ��9�d�L�ʘۥ<3� ����|e���5��n
V~$��͹!�b
@ Tߌ�\�'c���%On
V~$�i1n�6P��4,�Q����W��'�)�Բcf�x�HZ�, ���q3HL�1p/-��}-���NHRxF� lƔ��M�c����#XN�w��o2�n�����9$[{^��o|����"X��[����fb�W�6?��c�!{p85/Q����ߝ��v�Y/�ܜ�������#oM.�����a�x���,����)>B:�Z�m�۶<��%��������O%W���c*����b��v����a�����pP�h�Qf�Ϻ"t�Z;��6J���Qטg�u2=+쉀�z���q��k�a�x���,��ג������q%�����Ժ=���]�_M�<TC���qyJT��rW��]��C ����X8��8���/���K�����aٔ^?�j�>���/���k���cSS�b�E�0#�4j�T�\ ��, ���q3HL�1p/-��}-���NH�}w"�5 �Ac�N�AO%^�p�c�g��U-�e��pʆ�)�x�.#P�j2E�?�5ߧE4��>je`��@d:�����{~Ϻ"t�Z;��6J���Qטg�u2=+쉀�z�蒎�Jy<��M'�b�	�)�.�i��q3\��L�1p/-����n��I�8z�X
3kZ��5ߧE4�핮�0`K%Z�Jd!IG��51�X�c�rs�i�����fb�	�)�.�i����m�qv[����32��4� *����|QR����c8?-+eNy���@�KT۳�͕��Y���:؁��_L� "mJG��4JQ5��fյ��a-6�Da�`��t����@|�)��8���e���a-6�Da���н�!]0{ɽ����c�������aٔ^?�����zyNc1s�B�~�%���0�o���x ���b��v����a��2��#��w,��K�$�s�Ec�5*�'�)�Բcf�x�HZ�S]�*
�]v1�_ُò������?O�y	�?�\�
-�#P�j2E�?��˓#��͑i1n�6P��4,�Q����W��'�)�Բcf�x�HZ�, ���q3HL�1p/-��}-���NHRxF� l�f~,q����#XN�w��oֺܜ^ۥ�W�6?��c�!{p85�ɮ��؝�b�Bϱ���,��ג������q%�����Ժ=���]�J�1��씑�:��KY�[b%Ɨ����н�!]0{ɽ����c�������aٔ^?�����zyN#P�j2E�? �X��E=r5J�Ӝ$����b�Bϱ���2�b=��_���x�p�-a�D͢q��`�L��F\�l&�c%=�)�]�!��	Ǹ�y85��C�%����ۯ�����Z��/��\�w�0i%(ξv�釰 �X��E=r�����Z*V�M��nD#k�˟ܒ�o|k�LbfF�5.]��۪	�}a�IX0F�Mұ�*ȣ����W�`�f�cKݸ){�"��}����@����p+����g�I��e�2�=Y��>{�i�C��-�RfJ�J|[��alD�� {Z���ڨ|����.�e��U4��\��P�%�+ Ixcw���Z�����S��C����B)|D/[f^���;��c���X K�D��t䃦�=���>��ڷ�y؛�"�'����"O��1h>E}#���Z��E{'��p���qU��r|]��� a⣃_BO������k:͋��C8�oFJ�u�S�c�7�i�2�L���)�J�I�)�z�����]���I����+��C#�K�"a��ُ�S���v�?�����s�cki`:Gu{�F�ï�y'Ƶ�s��n��I�8�}w"�5O7}�»p�[k����Cҷ��e̷_��yC��S8�k��m�ݧ^ �H�� iJa��������ܖAA/���G��=�Ӌ��rW��]<���,Y#A� ^M'��k/��m#I�A�5���ò����{��|M1�9$[{^��o|�Ψg��U-�e"�A��"�Y�{'%s�.W�jb�ԡ*
T��Õ���PLJ�/���k���cSS�b�E�0#�4j�T�\ ��ه� �4�< ]7|W��*��fR�9f2Pih{];D�yl��m��'A>�NjX�U�6j�"Hs�󌘓S/�3�	����;;��M2��<LC9s��� �*$��x�9��_ڟr��GP���*�N�^���\�}����� ��$A"u��p$(���%����H���=磡��{��1Y�[�2(���($�|�*��=| �����a��Y� ��|����:�����r����TH�_��^��{��|M1�9$[{^��$t�3��T�\ �͊�51�X�c�rs�i�o������
E$���K��U>�f&��'!msR������K�=p�-�	�}w"�5O7}�»�E�0#�4j�T�\ ��ه� �4�<��,����)>B:�Z�m�۶<��%����ZQDu����-�Vb� �Z鎬�������(���T��}���9G3;�hs�{�"��}n�m!t%qa(􆿳��@�A��F1�	�A
�)�𭅐t��PЕ���PLJ�c8?-+eNy���@�K����,�ǰL�[��V�1���q�Nv�iL�D�"��^�Ǔ�v�����������n��U�;��c���XF?;��`9���p+��V�)Ė�P�H�U�B҄V$�qn(�>�{��D ΅R<������O�u �N^Z��X]w�)��Tf��뻣[����7.�O����좺O7}�»eD��+÷ �*$�8�RX7��x��0����}%���f�㏨h�(K�y��!�$��p���BBNn�j�;��c���X��j@4s�,�]�G�`<����P.A�T�g�v���>�֔�n)Pf�� '���Xw�j�7������⪂!�Jv�tH�����vW}-�п� W��$0���>���˰��0������:UkG3;�hs���p+��v W���}q�!D�t
���"X��[��h�C��hA�T�g�v�i��Z��� ��WnAEP�n�o���5"�Y�[a����.t�*G�pC��Vܟ=�a���X�Rށ̶���Y���\�!W��M<�<�.H���{&q4-�+"4m��r!���.!T@>$��M�0���j�>���/���k���cSS�b�p�[k����Cҷ��e̷_��yC��S8�k��m�ݧ�G�y����k�)�;�,�m�۶<��%��������O%WJB8�^C
��p��*
{+Y���>�[6: �|J��q�}��k�)�;�,�m�۶<��%����'�]C~�̄��v���&�?���B�+�V�p�nB�W��`6j�"Hs��6X�:��p]�g3��Dd-�ʹ���?0K,�o��G,8}FC��>�[�$�E�#s�57�<" ���h�[z�WD$�GLq��K\�8�/ivڴ�tG��D��;��dPi���{0��d#E9�����x�C���|�cG���wn��j�M��D��Z?�G��	�S��-��U��?�d���&��5Zbz�Z�f�x�HZ��,e"75�EZ��s��rN��t"O]��!���c�A�L'@fU�X?0I"�`�it�M��f�֝_�j�0=N;]%z���5��Z"�'��G�<���,Y#A	u�e�2�?�m�۶�so����O7}�»�QNȮ���k/��m#�J'�!���=�@q��u���"6ޭ<:�&.am� W�����H��6�Br���N%'tF��;���R��C� �Y��#_1�|.�~� �����$�\՛��2�k�S�{ �d�*��M�,4#�rQ��G�t>��Kò����{��|M1�9$[{^��o|����"X��[�-�Vb� �G/�'8k�{��|M1�9$[{^��o|����"X��[�w�����3�/!����`P�0M|b9@��P��9G3;�hs�{�"��}k�����#�B���BD��?���gMsC�|��dkw�Y�z{�P�++�hW�w��fDu���:.�H����,�ǰ�!B�������}|X���zM{��_�/R{-z�}h}�L00:;��|B��J�#�pV��>.�3x�В&=�y�q}��"�"������x�l��1�U� �1�}�W7��c�r��]n��-��AmY�f���e����+��A/|!�`�(i3�tt"���O?�R��n���L�����+J���5���Adu���h;e��w���U���~��yXpo�h0�h�#"
s���
��y^Ii� 9Km!Қ�6��,�ݜt��ϭ!7y�x�ݡs�����m>>*��H��b��|fa��
e�3+{�i�m�T����q��cy9k�\,����\��ʩa�扈��n�T����j�>���c8?-+eN�CyW�f�t�1�M]�'Ƶ�sס�Wd�#��9�,e"75�E��W��_�ړ8���/���锴�;��|B��1��V�����m��g���*�ܙG��	�S��-��U��?�d���&�	�Ao�'�Cr�%��^�}� u��O���#Q�(o�rݧ���������ۍ@qAnA�j\�/���B�wj$g�X;p`��/���k���cSS�b���$�o��X{yAuޞ�����i���a�����Օ��qvdЧ^{�j ���X!�4V�H�%p"��RfC` ��\U9����u��B�bq��2*Q=F�k�mD#V��[��"|�W������Ϧ^c!�6 �ef�/EI���ā4@Q�/�`u_=3O�̃苇��Fe�.��=")r���ꀍ�˺�Q�����+�+:��M���ʦ�<��K_�0ß\iygҟ�%ў׫�Jd!IGG3;�hs�{�"��}n�m!t%qa(􆿳�E�� ��M��u��%��d�)bUB�an�~#&�rW��]��C ����X8��8���/���锴�;��|B4Ǜ,�3��r�qU� e'�ZX^�O�<�V�QK�}��"��R �@B	���w�|��@���� G�� �1G�끺���SD(�
��G��	�S��-��U��?�d���&��}����MB	����ߝ��v�Y/�ܜ���}��9��z���FY�g��U-�e�c8?-+eN;�\��	�8���SY�N iJa��������ܖAA/���G����aU�D�mD�VOR�)���$~�ߝ��v�Y/�ܜ�������#oM������c�����M�~��4e62A�I����Oݷ �*$�8�RX7���#g�k��9����4`Shz���{�"��}n�m!t%q�GWV`��rp��z���m�OQn��m��'A>"RX���N�[��|������hM��1o�l�P�_��� �Ac�N�A}�Q����G3;�hs�{�"��}n�m!t%qa(􆿳��	�,זz�V��	��y���˷�f�b E���6j�"Hs0�1�e��M��a+g�% f���ìq�8�T�����P�%�+ Ixcw���Z��[�nU��H��<�C_�,���� �Ac�N�A Ҳ́p��xkx U�_@է��c���ĽNl%��?�d���&�7�䧅��m?��~]l�*`Dg�8�Hk��|��m�d�6���!�=�ߝ��vԶ�$(�������#oMT�K�^d��+?B�OA{?`���v1�ߝ��vԶ�$(�������#oM�������G�Ȧj�E��g�Hb�=A�z����gשP5}-�п� W��$0���>����i7A�r����/���k���cSS�b�l2�_�V��T�\ �ͭ��t��PЕ���PLJ�/���k���cSS�b�l2�_�V��T�\ ��e�P�HPM&�*�� lM|�"D^���\�}e�k����b}-�п� W��$0���>���ˤ3��g��c8?-+eN�CyW�f�trN��t"O]�E�VmM��}-�п� W��$0���>���ˊ%[��#'�,e"75�E��W��_�ړ8���/��ݾ-/�;��|B��5\tBO��G�Ȧj�Q�ͼ���݁D�n��\��c���Ņ]g��3<۳��@�>�F:T3u��U��)���Pa�L����N����w�b�i�j� ���Abs��2[�a��o���S�cA��(�����H�Z��+C�>��r?j��h}�L00:o���wu6�_��M���!�'��أͽgF"?{�"��}-ֹj~bЉ�؈a�����1�R��j}�C���&��vt�*��]�3�@Dx?I�{_8�Y��=�}�VݨK���L����6�<Z)��;^�|����~���i�x��M�j�l܎#�o�h�d��JXl'�T��~��?u��C@�q2'��8�Yu��"Όd)���l�#g���D5�|��7�OT�,{�"��}?�E��!
O�k��S\���������w)���r?j��h}�L00:�?��]��J	ъ)��֝_�j�0=N;]%z���5��Z"!�%2��N�E��۳H?��~]l�*`Dg�8�Hk��|��m�d�6���:Vg��Iقgt��ufb��K���L����6�<Z)��o�B���/X*F��c�D&����\��H��$�)�vx�&�l�/��+�7�����n��C��ip