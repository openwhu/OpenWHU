��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�s8�R�	�}����pn�R��}"6�l�:���;�g؞U���T��ײ2��>���^k�/7�?1�(�c��ߘ�]���<�j�C��`��L&`^����8��U�Z봣��D��L���_�L�3��0I}.�ANMs����C^�cS���N�w	*D���y&�f��+K��[y��ڂS�O��6b\U����/lt�3� P�;��1�-��⫯g*P(�C#<�:z����uP!ߌ��˼�{�&��ѕ���jǎX������n�q5�(�+}c�)�Y¹w����HNx�IL���om�Q*���T�K��͛�����Ŧ�l�N�`�ě/:cї��������qV��6���d�e������2��zEI�Ý�M���A)a��4�D�h�1� ����;�Ӏ�md�L�aV���o�C��ɡgJ����f�P��_�v�h��`O��Ftl/�~8��Ș��<)4�H��vE-,b����Ǘ�Y����<�4�X#�Mwn��A@�r$�ȭ��J�w��<#�+�[�}��|A�Ww�=�d���Fz�!�`�(i3!�`�(i3�<VP�b� ��E����q�B�^��7ص��s�r�X�<\�t7��s���q��cW�sn�;��J8�����3(:�QuK͖!��x�	vy��s^�&���Fz�!�`�(i3!�`�(i3�=��W@y�]�� �OׁΫ3݁_��޲L�&�V�.Ю ��&\VI`,�ʺ�;[��+$�6ﳌl��t�1��꧄�c����E�zy�զ3�0�j,-�q�m��c��!�`�(i3!�`�(i3!�`�(i3 ?[n�:#G٪�t6�yG�?� }[�KO[2vj���B�N� ��b�FP&ׇӭ��!�`�(i3!�`�(i30R��=�El����W\0���JY���y�!��_��0_��hd�Z��N�T?wׇӭ��!�`�(i3!�`�(i3p=�n��ɬc��WN�����<�FxNߡ��IB��<W� g�[�ܰ0|]<w:���G]Fň��h��<�rE��"7HI�S�k�,�B���,���}0xs�Җ,G����Fz�!�`�(i3!�`�(i3tk��mrW^~D�n��������t��p�O%�+�}mIƾ�Nh�m ͠c�|�]���!�`�(i3!�`�(i3H������gf���)�:	<�J��I�s�(�ߜ1�*�Hg>pu�y�jI���뺨���!�`�(i3!�`�(i3�K�Ǔ�\=RJ��z��"��:V������(O#�e*L�E�w�̙	,N�y����~p�7��w��b��rH�>�S�6�0RD��}��b.�Y�PG�(d{��8ѭƦͯ\�Q~!�`�(i3!�`�(i3!�`�(i3L)+l��n�����<�fi
�׋���1�r�63#d�ׇӭ��!�`�(i3!�`�(i3�ݐYs�����'t-/�9D��}��b.�W�BV��(�ߜ1���ccnh?�!�`�(i3!�`�(i3rK.��=(M($FO�X�B�ei���s�61%=��+��>�6AcUgE�ϧ������c�$ׇӭ��!�`�(i3!�`�(i3T�[9�=D֦�ccnh?��sp���(�ߜ1�U`�V�٘��LТ��-������LB�����ɧ���~O�kQoZw�ןLYsȸ�"rR!�`�(i3!�`�(i3]��g��a�5~e��T���c��~$s�c��0ے���(q�� �0���h�)���Y䋇	���1��/z_�����h�[ѽ
�O���6��2�k4|��1+�l��r�����<�>�y&�E��}�y��X2��6Z)!�`�(i3!�`�(i3!�`�(i3ZHm>��.;��L�Oɬc��WN������J�A|������l"9�ۗ��!�`�(i3!�`�(i39�O��F�=,�m��B��sp���(�ߜ1���*ȑs��!��z��A����\�K�y؄@�!�`�(i3!�`�(i3��+�t2���zЊA}.��ccnh?��I,�D�y:#9�]�B�-����;���ԝ�i�Ҕr���7��Pgen�MS��5*��8��i�c�g���H�!�`�(i3!�`�(i3!�`�(i3��o��d<r	�%\*<B)363�8�.D�V�6�˅�ٓ� ˖%*����ֿ����Fz�!�`�(i3!�`�(i3}�E%|0�WJ�Slm�m��}����.HI{?a� ~>>ը܅%Gbغ���:�9��#2c/������=pds~��E&����Bsȸ�"rR!�`�(i3!�`�(i3c��N�wC����P�B�/.w�u�$f���܃n��]ȟ!�� !�`�(i3!�`�(i3!�`�(i3���C�RgҘ�I9�UC�*&�+�eؐ�����!��B���k�c��`�	U����f�7U�i�#!����P�>+�va��2u<�F�x��_���RQ�
�0��,��X!�`�(i3!�`�(i3!�`�(i3L�E��1I�OfUA`���B��ҙ����WH%���ܜ?n昼�2#:� c��(�U��;���-?}`�I��d`ȯ~��.S�M�#0NUD60L�(׌����Ƴ�����4=����f��b�+/ �M�p k
� �,�i!�����"��e����l�5}�
Z$��9�jw���9�ȭ��J�H�M ��,J�l�/�I5@�k{��� )<`w���'挒_�>c�?��ț�?� �عNUD60L��c�6�fSTh��\�ڰ���gLE�z�:
C=�!tC����ı��#d�F�[��m�O�h|���*c�M�B��; ,@�� T���,�� ����]P{�u�$f���SH��{?a� ~>>ը܅%Gb�}$��vk�,�ŭ�O�V2y/�q4T�An�� ���T�BQ���n�n|s�)>ΊՉ���6L�'�1Q��!7s�9��5�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�WOtl����m��c񃰮��^�3�Z>�=�G	�L�UGj��o��]v"5[�Gj��o��Y����6F$90�H1�����\��Hv��3t����k0e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���y�A�T�3Vl�� �̮��I�#<AuA1����v<<,� 2H����QkO|V"��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hͥ<#���vSB��n
HDW�Gj��o�l�����CGj��o��]v"5[�Gj��o�z^Fh&�ȕGj��o�R��(�.cGj��o��(���H�Gj��o�>�N�)-H2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�b#Ӡe��?�F��&k�ZV"���:��#tC������s�Q�_;�"l���c�a����9�ĒTC��0���M�<lbtsR�b�"oʭ��4>rS��w�>��S���Fl�p�7Z0D@X�,4�?nϦE�6���������;%J���v�_�Q[�1��*��!?9�~����p>{��`�'�X�څ�˺�ƒLX���!I/���r&��\���%-��]�O���.e��!��z����)P����(��jD!���5�Nn>��
�*�EB���a�i #�� ��&��*mm�!=�y����h�}y(;⟝*#>*��4DA�,#��e�o?�M��;]��,��K!�ۻ2�e�1�ΟÈ�bH\�a�����RL�a)r��fI����F�����o�E���^�½w�>��S�Y�)\��B���|��S��2�)�Ln|����O2qs��s�L�:�;�T?��{}��+�����v�ɢ/*0�(b�ԝ���ɨVu��7���	x]̷?��+*�7��Mv�9�I��P2g-W~���џ�_�v%䨉͞N	����V���
��G'�۰�����M�,А�r냸�~���c�6�fST�jf&�~�7���}~�N{`1Kqn���D���i����	x]�)�RV!�7��Mv�9�I��P2g`X�8�\џ�_�v%䨉͞N	����V���
��G'�۰�����M�,А�r냸�~���c�6�fST�jf&�~�7���}~�N{`1Kqn���D���i����	x]���Ec��$7��Mv�9b�L-���MƝb*��4�8�:r&@��j�2Mk�(�VU)��*��u3����r���B��jN���7�� ��߼
�d�8DJ� ��m�!=�y����h�}jh�6g���_�-ִ�fY��/��Sd,�ϱ��Hx�U����� B�&"�D���i����	x]�����O��}�$L�7��`6�^���g&����a������}���D�"t�G�8=e����wHmM>p��&k��������Ԗ��RL�a)3���ʉ����H7��jX�+[�d�vԌz��S!�zg�Z�$e0���0��B�cN���	F�o�=�e �m�X������+�ct�ǈQ���\�4�s��{��]Q�TT	q��$��<�z5��J��eb�hW!'!7U�i�#!����P�>;�Ղ��G}Z��2�p��Oi�v���j�������JM�7")�E�'3H��[e)�p�R\��ꫜp&C����/B!,�G�;(�B�T0�z$�}���E6sC&�gG��Hc�e$���=M��8�w'��(�D�&�〨����cZ	�M2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc.�
͹U�~09h�i�Nq�{5��]�0�lK'���Xw����Q4?���ʢ\��|�����o�3t�	g�y�mq;����z��r���]��7ď%W�����k��d��&e�_�#�gWr���q P�^�&d�A|�1�:�Ω��]��
��rE���ƪ�(����D�I�?g�f{ì(Q[nS5H�j.F��%�	�r�e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcd��q�G�+��T���jB�Fg�Y씤`��p]�=�_ZQ�<^D�d�OJA�ٗ��J�y6�N�f����d���q����c��� �7ht��}j"�,�>E��ۦ� ~�p�'<�-Oɳ�%R�W"������i]��x�]�V��֪zw�&��Rb��Y�Wu.��+6v�������!�؟�r�Y�}94�h�'n�^0o`�U+�PAc��N�w�Q^�MY:��Ok��@zL͊�q���1m��d+0�l�R<�q��f�}��h�'f R�E����F��j��\w��0]��0�&�ͭ�h�O�0K��!�t�'���Xw�,bxqX�a���C154�EY�o\�{�o�j�",oMG~������[�]�!����M[��ǢyP��C��?9=����5e.��xu	�>��l%i�-�%t̓�@��Q�	4G0�TD��ό���.Ӂ��̰�!�ўC�k������
L'���Xw��E�d���%��ڃ�������]�!��	Ǹ�y85�C��H�����t�Z�f����8���D24N<I8����\.WS�UE^����`y������&��f!�`�(i3�]2�y�Z鎬����y��|�!�p�������.V&��B֥/~.)��3\�R�F*}�c}��uO��������	́߶`(r�M$�*|�(���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc@�����>P�2-i_\_��� �yz��$6�D��L���_�L�3��0I}.�?u����4�GO�Lw��ܴ"8;�W|�.Ҩ5�e`��9|�;�Ojz�ǐ
��4�%Z鎬������_�,�[/�cWM��`�������Q]� _ό���.�}�
�?��(R\֎u����}����d�٣��A�=���ѝ�ux�����E2�DZ��.��G��@�����U���ܜ?n昼�2#:�PW���[f܏����^�]�!��	Ǹ�y85�C��H����Q^�MY:�6���;b��g��U-�e,%�0g���[�=�5x�1����?���Y���o�E2�DZ����+�@�Vw߼
�dr��mnD�I=���O�rs�i�����Q��^#9�<-W`������a�"Z鎬�������(��`UNP� ��b�FP&(����/�7jݭ�F���%,�������;���EWr��U�L��Z�]�!��	Ǹ�y85�C��H����Q^�MY:t�vd�T��T�\ ��yO�E���%�;���EWr�A����[�]�!��	Ǹ�y85����u|#9������8-|�D��=�g�+��[�V�ᑄ��Q����Y���tz� �U�
{�~j Ɗ�S�<ƍ]X+Iq��ݓ�W�����\�9�<1ݠ�m��/�v�@����b�z'hۉ)��d�7�qĵݓ�W����/顰�ݠ�m��/�
cFI_[�x���b�ʁ���Mյ�D��5�G}�L?��:�wǹ](UyT�z�D�RG�&ց�*����@Y�h�6�q�� O��e��8���&�(*�O�q�N�;r����2N�3u�HW��,��}Dq�f��x�����|�����j�/T�<�_K��p�ݚ�Н�(aw)�D���Z���{�u1H3�D6�ؿC�1!�`�(i3t�Ϝ��;9��������$t���b��FҼ���6��/�����:j�D�mu�#��bE�������W�{9�ݓ�W���]��`��[ݠ�m��/�p�c�Z�x���b�ʁ���Mյ��Kx��L?��:���7�3mT�z�D�RG�&ց�*村����n�h�6�q��~��.�`�8���&�(*�O�q=#{#6����2N�3u�H���;sY��}Dq�f��x�����VĽ.��NOj�/T�<�_h~5��	<��ݚ�Н�^	O\�)+���Z���{�u1H3�ke�"`g�*!�`�(i3�S�%~�H¿�������$t���f�A��m��6��V(pyL0D�e�qT�e0q|���/?�-��r�IHN��R���
�Ŏ��Jo���j�����7�<���Ŝ��^/���lQ����Y� 8�*x&�˝Sz��E�4.@�^�Ɛ\倲��y��lDQ�4��c	��Ј��9�y��Uv�ݚ�Н�(����/�7!�`�(i3!�`�(i3!�`�(i3��xAE�g��Z��\_�!k�,��˝Sz��E�4.@� �o�X�l�i�<�9�/��K���6R��*Qݿ����`�|�XCtKN��ق7�v�ԯ��Q[R�7�	��x��ݚ�Н�-�;S5b	g9��7^y�,0=]^	�&J��ס#T�&�K'm=�;b�-�2��;�P�t�5���W0�]��e|)0����)�x���3�}@H�[�{�G_TT7���1�; �L�q�t�MyފVZ鎬�������(���f���k�,��cEp	���>P�2-i_q?�y��`p�~(�M0uѺ��-�ۢ	:j�5irAz.lY;�e�O�!�ўC�k����}o�`�����<Z��u�=>&S�XQ�� ��&�>&S�XQ���A���Q8�w5+�uh����M��혅vº��żפ	�?9Pjp��17e��:r����ZqJ?�d���&�[��N��h����M�&uL��t��B���N�gl��ܬa(􆿳�OO����˝Sz��E�4.@�5�J�_C�E2�DZ��j���R�oV�.�g3Zv���� E��BLV�^fkӂ�>�GU����,����#Y��9R��<��������ޝ��Jj�C��5)w�	����=2�L-�$��^)B�!�`�(i3�E����Fxy0�u��?�;���]�Y���v�岦�%I^:��%9&���;���EWrqi}�Еi!�`�(i3��os�z���+x�r�s�*�I�'���Xw�f70���6Q+�M�2N��n����eT���_L�L���\�7],)�\U~܎VV���~�26��\Ϥ��R��!�`�(i3�����5	�3C���_����$�Qu�HZ�;֐��F)t��1�E����F7�PɆ�˝Sz��E�4.@���>�֔����{��~�26��\d??�A��?��s��Z����+�J��*`4��֡���A}:h:
���9
!�˝Sz��E�4.@���^Ԟl=�4���܂}E�$5��յ[+8�`��CYތ�;�0�s�{1?�a�ؠ��<a��;b�-�2�Ŗ�	�&���|e"V	��V}>�O���(Cq_c�!
�T�r�5�yo���_$�D���|���޾o;�fu��r��R�͢��n-/�)�=� �s		̰���a�~9��tf��!�3$�J�5'!�`�(i3=aUh�����}��!�`�(i3~�`cC�4�cOF�{����rs�i��:5A��p��0�&�ͭ�h�O�0o\�2���ϵb��h�1j̲����G���y��lD���|�D+�G_"�|�2�ݚ�Н��]��/ݐ=k_0�b�Y�{'%suE9�+�偘�̰�!w���B}�4�N��<�s�������5�*M�yλ������ݚ�Н����W��Ȑ��?����2�7G��������a�~9��tf��!Z鎬�������$��'ѧۢ�%N_PS�^����d����B��ϵb��h�1j̲�2���hs���I�WEĺ_A9T�7��q�4���=�,D��O	xc_�q�����\��fh����G �U�'1�"#S�K�.�� ͷ�	����x�{���:=����a�~9��tf��!Z鎬�������$���l�^!��'(���4�N��<�s�������5�*M�yλ������ݚ�Н����W��ȐQ�rG�LN�ݚ�Н��]��/ݐ=k_0�b�Y�{'%suE9�+�偘�̰�!`�����B����t��ϵb��h�1j̲����G���y��lD\u���Mh��������5�����}Yms��/�u���4���O�>�k}�r�,0=]^	�&��|�B�����Yk����Q�Y�<���%���!X�I�Y;�jmT�#SDn��r�Y�B�{�mo�.�� 낢Rb��Y�WA���V?� h�ҩΗ/��@����*��Sx��1SX� �uE9�+��!�`�(i3:�HCaIMl*h~U�?u��!���c�A�L'M�M˫ɒ�2'�m>v��v�K��������ȓ=�^݊��}Dq�f��߆�p�h��=�64�+�E��&"ʞ�^�����t X��ݚ�Н�.��J�޺��:p~	���; hT�!�6�ݚ�Н��� л�qe��㎊j���Ű_
��m���c�A�L'�
nЯ�O��wӨj]h�O�M:R	� �}�휨�:����D<��5�2ԗ0z�cUL��A��G� ׿`HڛuE9�+��՝� s�#jE9>н���U'���>
A��%��WG���;� h�ҩΗ/��@����*��Sx�]2��,� �޾�Þ!�`�(i3��n>�ϸ��r2�C��8Nԩ#�8� &9x!�`�(i3�����VVw�⽒�����n,��'�\�n��*��[�ݚ�Н�����l��y<��`��ï��4s[�';��#j�ݚ�Н�!�`�(i3套�qD0�d�i��?+�Ɩ�������|e"!�`�(i3��jVѭ@!�`�(i3�2��}��E2�DZ���3e\�n��뾦�!�`�(i3���%>�rGO�D mWN!�`�(i3�u��A�0�Ή*��a��2S����R�	��x��ݚ�Н�N�D��泵UPal�����_�n�֨ƜR19��ﭸ�2���5��03���$73�!	�Ø�e�!�`�(i3��Ě�����}Dq�f��u��A�0���򴶽!`���*1$f��_Ub�F�S�1 ���jVѭ@4���kc9.�}.��]�E�i�m}6O�D mWN��m�5h1��e�?gm�#���T�s��R7��i8�
���]6\�4�@ �i5�Di֖�߾����k$ �/ٗ+���H6)�B�K�N
�����7��h���,��
��+Zչ�߸��S�Ȍ'�� ��@O�}�,%\��w�T� �f&���#��uގF1h��r��`�@2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc*?��J((