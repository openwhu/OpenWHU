��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω��U��}��x�� �� ������[���a�8%`��4�s�6�XAoeu��a@����þ�V��1�Wqlw��9�K���m��+o���sp%��X�����b1Ø^���#K���lӧIA�a�V��R��tv�Τ�䎎��J�'�دv)h�V~�$v�p��"}�v\-8�������>�`)���a��rl�ʩ{�Bfळ��)���X�$� ���jǎX������n�q��}�p� �Ñ�]�*�p�㈍x�!����Y�f��a�Z��Vb$���N[E�=����tL��	Z�G�a}CK�fC���4�O�"�F�È���_�O��<$e|����w'��1�:�Ω��U��}��x�� �� ���������	x]̢/����wЯ�mڍ'T����X�w{������:�%�+T%2q򋙔�M-US-�8<�n�У�Ǝ!�ѠV�>!�/�7��u���nEA��0
!G]nt��⫓���RL�a)'r�Ӟh� Bg�3���M Ce=6�([a�EF��7C��Hwɶ R�p��4�s4�o�qR��p������M<D�7�s)	w�N\`�a���!4d���-sk �0%̄sb�� bL�k>F�泂�0�V�@���RL�a)�G{�<��mߍu�M9ts{z>�z����H��~�7C��H!�������0�"���L�M�=o����"���	x]̂�FQ�Nc�J�M=O�A�+�4�Ҥc���8�:r&@9����DUɐ����D��)/�F�5R�yב?
~}�k�������E'����)cڸR��wk)4�
�u��w)�S�3k:�(�-c�J�M=�O��yt�C|�jw��[�8�:r&@mj�,CϷ#�߀�Y)`�k�8���҆�|n���:�o�E��Uu-M�rt�d{��}lJ�Й�m��?�Vޱ������{����VjrHS�w�MH��j���r���+W��YJt�,�y"r� J&g~���c*& z�s�ђ�B�~f��0(�/��$ }2����T���Q���!i��ӯ�02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vce��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�׍E�+��
���*,f$�7Q0- ��Ck�fÜ�2/���}����сsU%���n��/���Û�E�tw:g+��T��d^��_|��3g�ݜ��s8[Z�`
5��*�z�������D���J7"$�zV���a�ѬL�1m��+Y#_WӇ�s8[ZΑ� �}E+�6�L�r���{b�2"���Bpш�#w��q�©���B���������'Sea�8���`<4}��(����5�2���[@%����nEA��ȐTo��qNA��d��1�:�Ω��
�/�r��]���P��`�.�D���J7"$�zV���a�aC�h�>�N{a�9O��Yk"1/o���sp%r�M$�*�()�z�������S��"���[��ҋI7��-5�B�wj$g�b9���1��]2��2�F�PY~�y�����[�JHn��z���G7���� �����x?����k�c��`��'n�^0op40�zɈ�P�i2s�4<��!I���1��ݥ�U� ���_
`[~&�x/���i� � �	{����0�&�ͭ��|g�Y�'���Xw�f�VHF��>BH<M�z��]���>����CΫa��������-��%Mό���.�DsQ�V�r[%�/��{l�f|�ό���.�q�\E��0�X��?��Z鎬�������(���`$�P.eE���lC��U�T�\ ���A�������Y�r��@IE�U����S8��Ѽm����x?������lC��U�T�\ ��Tǯ�!�tӱ1R�m��+e�(���n�JŬ+�
���<�s9��0�S�&�����"m�K7{�>P�2-i_���F�� �yz��$6ea�8����U��}�o���#V�2�Ў��}�
�?�����}���=�?I��)^�q�bx?������lC��U�T�\ ��i3�|)sՀ�T:���V�s��ҟ�s�_E��V�no#��٠R�^Ƒ����"X��[��Q[R�7����n9�yE,~��7s�9���o��S8��Ѽm����x?������lC��U�T�\ ���>�����+�@��ZZ¥���5.>�W��*(��F���5�L�1p/-��P �R�)R7x?���Ա��E���2W���R0�����wc�!{p85c1s�B�~�yӮ�)��	n�1tnzʘۥ<3�\"H��E��F*�L��!�`�(i3�2��}��+�n�)����%�!'G�+R���o��_�Rv�䩲$����x|e�Fd�G}%�ȏ�%|������"sS<�0�zG��� ߛ��u�����j�Bp��vdN�<@Iv��nt=:�v��؄aX���$���͜P_�_S:g�RMm�o��'����d����3�H�����Yu��� ߛ��usȸ�"rR�+?B�OA&k@C�Ɨ0z�cULb���H��u:/�ˇׇӭ�����F��O���uZL��\z>�L���$H��)��os�鮊W;§`����;8Qܓ<bm��+�Z����y�����=pt�iZ]XF�hx��G��N����p$��<
DN͗&8�,�fC` ��\U����z~��5Z����.��֞�������i���a�����Օ��qvdЧ^{�jf�?ǉ�=^P��:w0I� X�1�8!�w� �O�z���Ԝ93����gh�䊉��	��J�6p�N��2��,Wc��I�W�"�Ů7�6��,�ݜt��ϑ_�������� "5�]3Lv	̅���X;p`�(�������0�&�ͭ�U젩`#�4>?� �1%��C����\P�ʊQ:��IK��<��_(x��`g�%Y��̗0z�cULb���H�i�'�/=n�t�{#	�x����dЕpב�B��P�C$ �lTN��I��!���c�A�L'k��< �A�f�QF 2VU�簦!N�'�y�G